--This example file is for demonstration purpose only. Users must not use this keyfile to encrypt their sources. 
--It is strongly recommonded that users create their own key file to use for encrypting their sources. 
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
pqJUsYqRafhpXYLZUuCnGKTR1Y3bAa/VH2fzFuOGdIkypFSrTjsANM90k8iLD+UXl/IjnE1cFqAl
Wkad3CT4WyG9Zl2MUmwAkYzVp77ivJwH4XQOHo3ZtrNTfhWkP9bOQURwfXsEHWN6osLekfr6MKR0
lOoSx8jcmMjBps02OdA5IfA6Tfb1mRJSmJ9pQXsEhGvxdcperjEdE9fvWzUPnuCOP03wlOuWop7U
iNydOu21p0e7lLi11hcaW0YhCRqEDXh1Lrmw+QQvrXAWLQxOY0QOqBX2wPkWcp2DoTmdwbZu+LTy
o2IjkGTEB2DiMOHrbUXG+RjRAhKfM2dO+/MMrQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="hCSqkFgvNn5+ruCKU6cQHR7rjr2psfqzeom6VZkUmDY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35504)
`protect data_block
JLfmQzf2mRB+jzdGC6ZM8sTcR8IhIwJSEvrfiKhZt1eCdtgVFf+O5v92kCtawHRJMPc4r86oqiwB
q5vbFSen8i3YGMgqlkitOGu8oLaH0jZnTt4VMusfMcYAGNBkuv53OyKxkJluBYs42CVIeZCuIyUF
YwA78kaR+fjjUtsX/CBSAoLcK/FNw00YksF3ZURWm0FxgiEPd6k0bfRmzcqdPF1klIac7juRpp/U
Wfkq9GYZ7dx+VoFwkBnn/a26nzy8SmEIHjErrbHyddePXo8TFojW//zPJ6MaH5BaWJsg1PXuAuKH
vp8FV0P7rC4qDSU38N4ZgB08ldimTP17YR+XRBAEZhZusywCfQ+oL1L3IUAk63LQB1wu8B08X55V
oxTctdIFRtO52BbPQ4O65NkrWHXZRoCginDEIRs0YTS079D84vd+kx836P9QLBr8ZHJRudelD7bW
G6hvuE8lq9nIrtnELV24S71XGW03wR5YL4T0z8frxX7zKKxBcce7NKyUnPfT+JQZvlA5RYMNDDF/
AmS2KyvY058tGEZFLj0knLh79N2a5msYOw3zfNYV7KNqdmfapC45shw5psUbMxFeJeFBMw2do6DK
PpChF4R3QOQ2+QEucxXbAlDCOQpdnSYeK6/YmnUbGJxlDMhNxfHbntijkuBEyBW4eOJ75cR3QW0T
CiQjlQmlDebuq7aQgedWiBe1j/Hs44xIS2ZjpYL+fAh6AR1F+L3770rrKd1uA4Q+q7yeh/qsQoxj
Fo8mzBGtKLVQEojito5VSF2QyaLtS+wi3DXvXYl+BTafO86JHxwBl8iIp40oe3BnL1Iy7b0dx+do
ueQ88JiMpX3/qVO+GRidVO/EYm6NA2d4PkWcWeJUj1vh+T3Xtj8oV9/2sqfPYnHYir+ksTYEJAiB
1PtFxyr1OyLqrZPlGhWLXPJmUkfK0MG3a74RlFf/j5D+0/W8iM0+/1HN/a3lFc0+LoqAILx134Hj
3eSj6u2vuIjpLj2ac89D2TfvAbFU26Fowy90dSFy6N0TbHLmJkirV+IqiW/ywdhpwtpJlxXpOSLc
rEe6LL09dpcPf1GTDjhw2IWEymcw8jD3QdBy7rlrDuu+PI0ApQIXhFrJbQNrHMUrjvvSyS5V7kuC
5JcmMU44ArkCpJFUrOYDQXq1vQ5PFCjkokIIzjCXHUWRqfW200McwmoUQOG7Y8rd23KVGIu+50+F
4+IYqbfHnTUVLpuyapyxGt7Da/2XV8fkbxoUYwvNGR7BsA4Aeik+v3J3rdN3F6GGhJDd5r+d62fW
efMJkkMwlqPEdC0KrHCVwPvlmh+otBRS7sXhv9BYTpBRpuy/86qB3VuccHVCEs0Wk7bFj5ipvUi6
QjFIQYMlfKnJJ7ZIPvUTy19zq07raQYHWzyw42cJwbjYPAWgEx0uy8wI3bPaWwBWujkhN1oRfIIF
7vObB8oYH0zpf39v76hPuPe67DjqqIn2MblWMMGgWF8QX1v8ES7Wtedh8jXiz7ZpJwmU0vQzFU3E
DCulC8WoeyFI6DDqro7wDeKJGW1+LbqV6PAVuOQpk2Zzwsdh68uXVMjyUJOJSZQEd0iDg1WZc6T0
kMCAu7yE+tjO82iDPNHO7mV4J9klY1FLBi4eX8ZxPY7t73+TLa4sLcc2WRhjU1lB3aJudaBwYjlo
ajlE8uzXgcNBjMUMqx9c/r7RF/MtFeX64jWUPejrofXiauUD+mJ2W7qdmw2a2KN6dcgP+ZqQlPH5
FYcji4elwJaADMecc6A29hNHfgE23DKPfeuorxhsg6VHuO4WRjBLWaNv7u70K7Bo+S6AtgkFbSec
+SvqrIFd+WMY8ICxRBvSitF3prvuKULixQCa/wGl52FTiumiirX/fRjc7uE8T20Ux/kdl+d/9AzI
xeoU5dqQpEoxYzrKDUXBpCpv1AmvOrzSjJyZP3s52F1/rNeYFfkRNgTymuzJUY0mCBTANzW+wJfG
+vqH8G2Bl5NabdGXB1Nk1xODtS1aMhCYJxBtzVq0LiBqECuUNeLNl31Leqg7LyLMkxFrunGFsypT
rFqP7TTdl4vrTe8vBA7VqsN8nN7zDjJtpKeZtlZBVXgcb4M+pTnsSZGotKZljFtAUqr6DLEsc10i
bNsUZps8lqFpOERK8VYl/VMi2nRy63nhhWgLk9moMOc5eEmnnNWoORHZbHhWurdtgYLZgsDiiDyh
G+mLizYcUC8BiR+05yM5nVU+UdjcDTv9jljfJzW1vmXJ6Lon8BPDdTEyZycEi38a2JL/hnFhMWVT
HEtvfaPLG415c6XG0mnHg7BXZREGwh4oNv+pFEN71j/fEHtUJiH7aB3tKJxNzIcJZwcsbmCvzkH9
TNrnmAeLa5ADKrLfn5uMW7hBaKvOJDKLTjAVue3gxtXMSspRnVP1JM/Pi0fcs2gnIuE9i8YW+xZU
F3S9UBik1oIwCostPcu5R9guhrdU5iuR9TDhlitsZM4zeyRyFYB6bIEjoGKbNyY5+iHhFhV5CV3x
/MfeEsmrwyMRwqhfLAQFNTeBk06A7i7eZ1J0qPama+YZBB6tlh5BOTKeyT9Y9dROaXpG/bqd6KPK
mB6xbaZUrZjXRs4u5USRIHeovLeGWfxZx9OAT6aZ8KbWuKKzfbZAWep+I41sWB1jQsOMaV9IUucS
TbuU1Kofnor8UtHOAYYUxjwwXgP4Mzlqwp+qdqYBDAU4u+WZafmybdcGLYSAAuNxogVqH9Nx1+Kv
6yFZTp/inn1/YDwSlB8h5NJMFy+ExLAO5mDSRTzy6hBTRfuXHflqB0dFo2rPeIMtWfJYsJS2O8F5
ms82okT9IMsi+d7ZIN9BZvTn4k+zSTbiRTQlszXJZbT18qCFy/FdlkJSz4lMBbUkRFFDpkTeGe2T
aVvOYJp8kF1a7PzsIA4Yvr+W4kNo7MIVITPXmQlFcmluFaS/gFVI6VQtrSrJ9T1jXGWZ0rBcm10l
FeXAqwf0Thm4PDaFXOfggGT2vF1eE460qSBtUYhPW5k0Sxu9zLsBFYtsWTo04eXKk79Ib4O+RP33
2iCMMyzavRZ2o1PV52eiPPS+t29Awmp2ALpM5qDBmnTQSNQOQgtBOyaBOm5hWTo/5s11VOBV5KVO
aqKZrRZpEFTphmHgaN4AMlYbRaSyUClwNLoFRTBOWSzNzuBtOKfgktCLcFqG/etGPv8RXEDKwlzp
9yGDum7U4/FfcI+78XNKOq+jW93gJC+tZlkumCdTOvrznR0mqfDgsuWsC/7+LWingDwU8YGMgO3O
1ffSQESLGtzBJfhMHt0d5M0V7lL2pVEwpzZXT0Efw8CxJ35MRO2qajHkTShN7fD3OS9KbEkJGNSl
JsUCBzJewwV8ulHINWIQ2nuUspwc6pWPlVYdf+e2fYoRsxe09Gf/LeB8NoSUJmX7NZOVfkQHCv1G
4/nFWeWc59oPMG770Tm0Dd9bghOEj0w6VuPYbFhRG2DtrIPDC5Whx9foXQraKaTXfx4fJNiE6DXo
l2xDnuwEcClKqZVlnG5sXCv/1K8agw08Z4elLEFfd5JtoowaVnChpFt4qOq2cpIkeBm59brzDfPB
jgODJRH3pnj2571SzYMTZsfNZpTWANZDZ9l7BAaLF2KJwwIFHPEsURZZejtm8Yc5712QMIVDVDc+
T1Ho19FxEKSJ+Lfmosm5xPAz+r1BseSQMzxftyyIzF58brTzRAr/oUXXfORX36ecdEgU3+sXkIE7
dw6pXcSlfCRAd/tCexnbTn/PoZpIkSDh/fEzPDv6rHVkj4NbPRNMHy77ShO7Moax09HsFvI7Tgea
LYo0Lv3LV06II7Mu6+u/iU9VQmY+Yr/Yz3lQAOYlBOK5prY/NIgDZFa7mPp0z7IxtBtq6ljKv6eI
ELRD2wTtKZP/yfIInjaw0UpPIUOVh6ketNkb6Zm444j3vsLdfr+e0Doyu6jz7mqYB+w+4J2tCuk9
KDYiEGKFwFr9F1omHIEy9y8d6VmaZSbcX2skOv6BEXuIvUdF4GNcCiXkJ7Xu6zV5WeuxpAvQzz/G
1gnpW65c6i7VDlDEKbTN5nZn/VgcX1eucquKajshQzCghaRxjCAY9QbBinXyb9xoqPmMvJEgFAGf
Hz9sDxuvqT2eFYt8ViM5QQ9qG7Ou4kRMYe0D6Qo8li+LKeBTCHamSbom8KXxMbXwYuJDYVFziLDK
Frs79cPlGrTizd20HPK1oTMXw3PFJbEyfqzaget2echGcxjliO4Zvh1UoA5IcN1U4miOoYoHBt3E
dJDGxO8xVYUVK8QP6qmmfNQ2OyWJYmyRC7C4pi3OIISy5UrrhkjTBGxdMUCT6o4t5Bcd4dQYVhjq
rIfJY190P75ROFfTx9QhiZff5yzn8lPjSS9k7OBt2I9tFNhD7iARXHErE8sdVCr3ij4tHcSVVzLL
t0N5BLk6Py3W9GQxQc+IxGB6PYIccoeMhA6pzmRFQWbuQOYGWZuK9KPv+r889YtFKdDcKYbuOind
kliTjATN26toYhE0nnCF23XqRGMyqMJ6zq4kg6AkeypSdD065HU9KIqYy9pmIbbIDqAQmLWR55+5
NnFoWKfEfFwkFHnDAyQWejR+Q6QASmtBSuTLNFxYyXaaPEMF33nuqMylnXJi95Ji3WUBQ6GyFywA
oBV7RGhUPuDMWv1L035buCKVO1XgAXPX8X6C92AqRq87ttDgrjicEINdMzfrRbDOqs9UlI4JOBPU
/D62Ny/rZr+CU2/GhIsyEkDWtdqIM9jMH7ZTxUuFdl1nK5MY1YnfFVmfDa9mRQ6+G8Ego57k/xDc
vzNFHOIzfUW7LL2bUW8VNX5QNfI4L2eoxse2w8Fw3kfPUFrNDj9Ra2QF/Ny02vUMWCl1d/sDmPSq
a9XcZosmsMox0h38G0ZCrqzUFvNAxaj6Y2bSoDpST4zUqwQyQqbNDcACyW1qHYy1X7mM8HBpSct4
/o+2XBA4qcJaOcRY/C8Lq2pUU7251TVMqD1ZIOWndWw3IY7NOknzfuTAmImVqZ6RMgm83TGESxkz
x7n7MSJknF2vJUil3xrh+V0tNipf78jh2/tYSDtTgdZqMMHFFtv5AcexoU8Gi48+k8zUIS+f/Dcb
lNxJGEQhdHL7fROQm/EChwMb6Rsy4WQL+fzKTnH90zJnRHdxox6Q9HgSmL647QAUSWCbHTkAJjwj
oP8y0+Pos6SKZgWu4Mp5Xb3JBkkTsCzkQt3BAxqptMeXsdj4DiCa7cBf2zyiKaBbRKa7IpKooK2h
Xf7wk3dpvOpFslYeFNFknVM4Nott8Hoxc20Y65LPNP1nQWa5qRikM+5qnGRPn/vWx1wPvMnAXEH0
4BfryHEPPB1UDKSvlJgM1iHWnBsQPBXfYf4WXaWxOs0lnJwzGiJDWaHxVx6qKBET6f+ED2gC9cSe
oiw55Y85fjJ2Y5/K4DgEWd4wsutJ6YHpSi83YkWpm4Wv2+Xt9u9c3xl0Nheo3lKlS4frfFK04jsE
DggR6rH5pdTBLM0U90tbzM4UNJ/lYALCQMZAWoXb3m4+PGe0AbqAbt4UXDZz9NlYyxhNvBH/s8Lx
Y0L6DPKLqJKSbVv2Ztehjz5JR495ns1E0bmxfa/o9xoqnNOu2MfQE64h0LhWVqIN0Wjb5BXRKGRY
l+UZX2/ONyJMcG7RWGWwYGKq3uBiXDipQsmyiR/uGVo8lSSu/D6qondhjJN9G3Kx1fIwEx5sC9o4
96eaBRqgBObHNzjBBGzcK1+StAZ/Qoh9gKMnwHi4wS3yPCdGTnTUASaGEW4823Ul9ZCecf1ro8b7
F9+I9FodWbKiVjKriddMhWZbHM1Ecd8ACU4flv5uyQ0J3K4rV90++M9JVjM3DNNJuHQv4BZH+mSb
aiYMcoSD8v3Xhl+x9DXrprZjDC3Mikd+Fb1e71Q+Aj9NpZYH+SGYg3oLa4wRdUVaEWEhGKGgvpnM
n0HjmoSMEI8MurET3O/iddO3Cz1bKPbdUfzTWn8LJgyJfUoE+Yu3jdpFIG6W2f2QgAwYetLIjqJH
NNuiO1hrv+sgZTmjpRz/3f8PNPqxiFceuD2nrSzyBQlpcSUqvdWu5Nb/AncnkPBtEfIzh0kRFV94
HACAAML76F/jH3Wm4L5AVmDWHS5wCUxl/qUjWMlvn/pofaaiNPZw4hmG3bP48yiiQKgXZ7hN8Hht
HbiucKCpN3L/8+oQVyDGQwwGCPhd/W9w+WgUEBMDLMv8ZDBcQWVUPfAoWgAjWYN9t/NKgrrZ3mHP
hG587LvsrzZc4LIOvnFx8/2KqDMZMzEU/9e9xpMEZfwEUi4OOngx4UeuvGeDCn7TLwvBByEjE93P
u5rYLw3udjDHBnLvOpKIwKi+aHdosL5gd5ARr6I77fi0yvEmw+lmSE9+T5LZI++o4LsU7LipiNJy
er7v8lRe2Y1G5sbaavao5WOwuqZqxqDwyWnInv4aHHEapI+ETQoJJH12VuIxygvirTTx9AAoi2DK
MKgTJjaAVCcGNGPI7X6sM1K0CU0DSKjQPKJwoTr3OQrC4WiuYO6tSorY2mMvUA2L18+qS7lXzATA
iAQq4AMhT6CiJ0to7idMRmicgWrlcbQRQwGDUjjGiG0QIlCfZSVS+ssj3nc9992sfINZNzHI6l0O
QEzn84C332t6RQfMHNotebKlsPQ8w5XkLtYrGxGiTXmx7NV3NtbymwQ7ImNl1CgQpVauAlZQs/Sg
a7BK0qUoVRYrq10l0yGlMs1NWkc8wAs8oQMXc4Yi6j4rnJeqQCBUbYVDMY+R4l9l6pUWItGrOaNX
G4EdyP+rpVteoa2Wq0VRaLrpy6++yyXjv3KMEEkQgQKbwILmLFGJIZpwdyzOxbU2ZYoSLPiuRX2K
8V0cM7Mxf17jXbUWu4wmBMLx3gnOSoS3Ivl6l8N+yV3cF0MsQQzQWobHgeL9MLxwdPGNsg/ovS9J
+Ql30tQ8Y8l8S2OaR664hlnGcynRLKHUpmDAiuOUWkBnvv/SE9I5ZimmY7mPqH9+k3nL9gOav6oL
BB2PqSywlrMiuIssyu+gn4YKb5WNhRTHE2P8u9SXMVSSPcjMqUz2qK5pgKG3ma8NGvMVQs8OzYqd
BDfBCj1HlXBuXn0YyNitEr9XyGVLrECuKtZZy9H/HsoME0tGgwnNtEyacv5cNjr5sElc7aX/a612
Eoj/k4uJHpaLgcxmmo2UsgB6NsmjnVfpO+ZbjOTIgWl8GKPVvyrBHowXqefia4eE27PfaIhjUQdJ
r7nSjWf1kjAM0gLZz/7loy8OBeoGvFBlVH6wkdxyvMeGzKbKRVvCz6ugI3IpeMIAXcdHRVhIV+yC
npbyClXg6vvCrEDNjz3arYrXa2FMBgRahPkqUJ9sPzpNtPyVmvNYE88xOZzK7oD5Xoy6WVKTcGbM
VHVpoHAndPbTx47dGxR0TLQcFHzudpuHShUD/l6u1wqbgcUbvS3a5kZtPcDdvIWry7iL1DY8d1l9
vn4tZqrU78BmFXw0TRUlE7DRlOuveVdblRmVe7Rc3kNcrzJe5DG9z0Pl8YtaMUl92H7RJci3hhWz
WQ4jtmRAhYQax0cgy4XpTjusghyD8soGlMqHDUGQskVHJOqlCfsB6TmqOLXmlAWuaBpMj0qoiAtQ
CCXXPJfMgqorP6HHmh42cSQqRYrSRJcz2hSp7Lmw6r8NG/U6oiDEnxwguzviz1Eq7Ey+Hb4UUlpL
cXpbk9lWAxx9lRkdFHd6clF4OPJ4aLDLHTLtSLFlUFY7LE+0+BsJGOK99VLAorw5Yym8j34GPRr2
5Z19epW5hURIBDVMyr40LSeiRlwBgfLFP6nfMqJLwwWCjgb36kFgC+HQY8FCl1StzUUAitSWGUUN
1UK1kxVaB4WE/m+x0XvuvV6h0FYlMUyE84Sv0b2myMzUu+UE9R32aREf9zilOiMYnwCwAnrAs+4n
D1pjEdf7bW3dvt1RpUUiSGvVsYH08REMGG/qx8ghcRQSsPeNB56I87ksg6+1IqnuyZXTroGiAfb4
XdqhuIGHg9SaeshJ3eqsnvE7A187VR7bPui0zWECuLTZflKlwV23Q9YUwUlBSabEno8lGd6O7saF
xywyOzCZWnQX8OFpVbmIDFRxftkxeIafx71bIdZ49Myo0wX0OAlBo6JK8/krETG5RQKiyh+dV6JV
eit9r4MpWAbACgmh9kByNJgAKsFjaUAGtGlhgefYAwivoKCCyw+F6s1N9CkUAKmoXrHHJbiJ0hss
6VxAWYXgt4UJdzV3KQ3lnpPr09rnMGJUQIsWZGQnMXJHKu4/uz6ljECH8r+AgfNDQVELLY5R11oD
GdnQusqz/oNrGjWpF1WfBuGXifhkPRj9WHzNsInEkqTvDbINd4nXbVlVgloo/3isnCpuXrEtCkj/
FGohG0FUhugqP4u9mLS5/Ny8fHFuruDeI5KSnEf7BmlF3sxHghLHc/ExlLoJ6fenKaavC0PzAdIw
AD96pWVtyblJq06B0WZkt+ZpAX3W/8wLVYZ3K65kD2fz/zc+HxbmpaabFeDg6KDzs2A3dLi9QO7w
HsR9AnbbFWhHJ+ctoKpchrCfqWm6xKzdhCyxO3GxWpCRIFWruqhpUnyHNeHcohwjfgiZquK+k+rw
pIr4sMXZiJYYRpaweoKhve8b/N1QEVkuiQDH/AG17lfFfWYPC40meu+h8tUeNqSRRLgmD8lRaSzx
9bhdetE0qfFbrUdJCdhPJvF7VwDAkKskJtmWOoMiWqkrZxLCfKm0VY4tTx9A3jyN4PAOA8935Wl2
XXnJGkBSn2aVOxpEPcz1YALqHPsuzkJEMzKvJ6a0HD6HNdF6HFT8M8ikU37C5mzDE9wCwRUi5spd
PNYJNf+wMvkXPVxfN0VoViDK9EGzCyKbs4D9no5PWqldDzh1eTPABwHQc6uIapv3issOGHkUagiq
PnnKGl6z8+xbAithwoFW28Ugj0QhiJtpFp1bC06Iyl/QeRJXkkZyJzzroRKi3gh/yULvu2l9Pyk2
PjBP5zB/vLVpb4ziv4AW3OKa0RqTYFqJnBXEB3FdKxcpxWac264B89wvehpTp2UQrfRPDVm8Q2/P
RcnIKg2QFhflyiI/j6xmnpTG7n7TzLUSQvVuzXtEoEJrQEs61MhxT2kaid9ys3iNQ6IFuYoTA9s7
1RLJ/AIvEtvEwDlaCDHHj/yczgUHKcEJxhIxvfJlHj9wS81jAJJgKW6kiIwuwqSkgUfFoDLM6z9F
dT5xjvYQGoPX1drt4qQKYAdZTMBMleqOoI6tu15liCwjR7tiMsT0zI/H7Yc+SM27IIJAFKOkBGzq
rTycIHdzFnHMwB6IMsdsXKtfeg+5dh/SAFh4+q9ec5KQXzpSeZbTuvqFrIiIV73GdBrNAv0AHvs8
jQsL1lyPTVFVIjTrDAHcCjSP5Qcbsv5C+Z6GpZdM24Mp8L2Sy72xqrdlagDKm3KvCtY8D/eHFhL6
OJDm85/vwp+M91QA1ELWTx6qAGL7hJsgGekcRBefldXpzkvswGLjPOuRleWBN9W9A4FW2hx5Rrux
NwMo6A3sLtIQd7ArKpO5ibqNrPKvusgtHaew2pA89wZlSCkMd5jQXTnBq9Osm+0HYNhMJPeDFybC
BygYjCRfwqokaVCL29LmRmgUVp22cCsl3/5v4HxxerSwzjrovRqO352Qi+YXKLDkREUcsjiMmA5z
To4k7to3129jDvDlVWDhQstiZYn/5XidQZyRTCMg1I9HBz8EtGPWPjiQ4HNZcKzDD6hD5sKSsYQi
Y7AJY3jzHevum9P28xLxw8xvZyNMxp9mhLkj6JGa2opb2qIuf0QPpaG4wFCyTISNkgMxWINc9ozP
Ny+G+3LAZsTZeCqSQM1oViyzBd//nEreEEJm+SCruIsrMFcrw9Z+JwAWKot8FPYY1IN/IgBw1wOw
rGj8cfaQHy7P2pOmE+jMkN0iWK9sUQzPdgdmSIu+ttoHWNZP11rbotCX965d/ET8qCsqVOWI4cHt
TE4fyzlfFvZ9IuiABSNwpCQ9lV1EMZP1Iy1iSt1to5zajFFuHL6+ujAyUvq8OJixaaD0RxPU+tnr
bMctL6N4wFPsOKXvRdiD3KmDeqMEQUmXe4Jf4PvaBqJysv/DWCpg0IAtnVKiS9Hd+kuuG711+aKY
fiwXdhmFpDSRdkHREcLmRIMWRnhwh3YYG1YsbEgvFJvadVwhZwXEqayf2kyRhGgpOv8+yls0v1vj
qGk4GWr9D7kHZvul7QniYBdiVzBB/+aG6xx5sszuOmgdbiPE+nwlUnqgQNq6AqmnRY9gNj/0VU7N
ZTsinY/T+eqF4w6wDaR9016ErK29xbdwcgmRVD8n3HDh6q//MQn1eT93HC9CcNx92Pt6pko2jB/a
QGdBf7TA08AAwb3B/UhwnRbaqd1efCxfS0ST9MnDlkKRz66vdBBtzyll7LV7AIPzi1UVPEOLRdvA
0Y6niHJC71g1PKpz1BmvyjSZp3zuVCNt1JT/0eIeHcKRZC7myRbLla0o74RCtQtjXmxIkMRqKC7e
xDtoe257KCZfeqRwAzT9Ynl3j+lqrkDmyv3NVd/fRyl44U+eBqnXRCvbSVma8BsXAkCW1SvGDsjH
N7PSsCU+PKodjRtzuYpuC6EyWvmcER0eAwNGj4E+WvpipHxgYPH+8Hf398EbylWKLnqVqC82Aqaa
RC7TRbXhqgZp/jAAvH07g5xOuF/rfXOVZYdMTUYsP+a3BK7myBtddI3VE6SgzfYFsnLymkaOJrGd
QJCV7iGRPcXhu7djevx7sZKQQBNa+5lkHKTn2x6ohR6/OkQJeuI4OUk1Y0HQgL64LGK1i1pUL/fq
OeveCDORz9pBxQ5PrHJYp46kAJPW6xFQkKVFeVWvS9CJE2LKdxH3QijOoWHj/bQsPtbqmV/GjqfZ
d0oF/0FrY542Dwn0J5aXg79zpW+F4OlN84uLJo8uF6wCDZ3vyluNNG2HUD/D0Wam2JLrjJ3I8x5H
ztrr6kJ+mFCV1tnG78AHC/NPT3uGm4wC8D5ulNwy1AavovPHLRA0GO6G4BlIy4B0f4VfYgVF1HY/
jOooPP2dTpj5a7/xjYFsmxPs/gTgV/MY/ZjDDRKhCSzDnehyzW78IBx7zWdm29OJ3X0JVNxJ45bV
9/Ru3cM+C3qEkccVjgZ8ndXV4Rk+Z0aUlJEvVTDDtzCcDh9XWfwAisjED8wlpfNHjNAWGRSiULqx
V45S9kiOFrTolMYe+fcmV+weKPUnAbkxJFwzbJiqjZjtwgppq01wDpOdjOCkmk5FILS7lOuGi7ia
FYC1fjGGV8JXdnvz3ZgZ5V7gJ1q5wkAcnEHmthU3vdFjBGJFLX1MocVplEm+jILwNUnkl8qkGBXh
VCpgDGjPFcf/mKxXiLHzO2jgZwCLlOnuhZmGQHSfMLRj9sLq+vkCzue64/cyrZzd8eTppv8zDlNB
cj59dFtyCaKwhr6jVKrq+Ya6wemGkX0SVmT924mM2OAXPaIormt70Uk9LW2B7KBc6UuJqUlMB5tp
PL1P6xnWZjeV0kqL7iahHMZ6XBPcmDyEwG0qlsOoXypvQhW+3Pwv3jPN6nGdlk3RP2l0bbvv0ozH
UJOyWwOwlsw2T3nNRw+DQJOWUygmaebk3Xey5gY+bbaPUettGMge/DO4BtvqllyucyQ0LXC7fs8Z
BL/za4Hx6Ov0VxzuetyYkAGvrY+cyTTeMgwa+pYxGw1QcH8JOCbWKJg431gvITDVb3kF7mrZ1GYW
v/fZ/8SSUoncsXBmc5U+qFg5da9p5hLvTFD15wm0McXrlyk7NlxnuY/NcyPOdpAXBJ1Ldb8fzs/W
iAD8DTI8HYcEnSYO3UtNLSJHHGgKjYed2OFhuDiLla0rrurtON9fC5BhlZuHtaaw/M43r77et7J7
g5zYYYc3T2r4bJvj4GLm+fJWS1wiIW6rTfely6ejiBTGzHiXVypMIw2JlT44DyZ3AhZfM2ip2OdJ
yj8zx/vg6oJkapf3Mvhnqngb3c2bmiA9F6LVK/3rOsrV0vwXnr6fHNqntVEGACoDGP3JFrGB3XAs
YmPmfbAcBWrsNjJdFhobgkwDMJOKKwUmS+/n6lXgaGedcgbRkxcS8jV/UgMZ9qaAAeUbALpO41CZ
M5Qic3Qm02Zsdq/WWA7SpKKBh9tw/FIsk92Jjk9w/5CI4zREEbd+eTjEcq2JbrzdwZKyuN+SLolj
VMZmiU8S1/xBih8DiOo/WYmDhxdiJ7HXF+4mcG6D+XOpUOEPBaoyB4c8pP3vtHIGU/98YsFG+zDN
RsIaGZXN9KimyDIdvccTAZ/yUs5+01xIdleJ6itUT2HzjTKh69MIhZjVz5tiISHVwN3NNnZWWULO
GDVOe/p1d9KXzGWonu0dJr1XuURGkXnXSoPr2iAJNFpUpJf2trB7hZkp3aEtbM97+ykaCby1jC1S
i2O8b9CJLZrJxvP1FPU0HyRnckxQ4xDEJ6xiiAWwlxJmANcPv7Gx9yJZ4ONZc69wFWKKZILP9YrL
dAJp0bSyCj1Wtwbl5uD21slMYpRikKCvB1nQk1LNe9ybrsRI8ZCMNqbAQ+dvH3PAMlkcsdSvdGv4
n0lov5e7URsmt920Fx83PBI+6X3O7/g9m3Tg+iAwZN4VDVLCu7frW+9YpFI8IB3Atm2xZawx2jtS
7L50h/RZDy9FN1Bh5YBGr9yQuDaTqRq/TENk0lnLp0OowGFVRnrrvOQeFIEQQ9IuKeJRmeEyT1TO
HgFhjm3RxCRXkqQ+Me8ZXdTHot2H2cp6KmLbQEUEnWzRW9RO870SEEjXRqYyOH7yByNJieze8yRE
IuZBBMbEKL/ypKCKUJvh5C638QOHfVTylM9nBvisdlU1MiaMQJFdmAOY1+VQFdQtIQpuOg8qRpUB
B7dJ3fTOQhxad2pC3HtNldXNddPQHOsGowpTqINgeMXwYO4cqRszJp2b0QjmGFha3sdbvoCdQt7h
tWRWlrzx1SWGUiFJgfA9EBqoQxeAPLKxOF5d1fqexy/5/1kS2BmJ1f3e6baoTCmg4KRMej2IIOb3
qm6yxgf+FHw0a3LaMA7sMCTqWR5pl95/aZDK1N8WLZYx+8hih7NU8DKEzTSjGVJwXt/ROxolkLQQ
ZNFwAx2TOua4W2IUjXaaV2NiZhZokRj7pMruFJEKr8qJp4MCbofzxPmC8Z3Zk2kjKyL1rRJKWaLw
95NhOe1mc7LHYWKd7JiFZw68v8N59mMC6RWpISnVAa2Pp50uZuJPwu/ixdvbqyuDbPaR4/QG91P5
uyWB9huq9u3laWJfdimZTkEOdF3WtLyiovXOH2l9UE4EEqig12pv1O5scqo8ms1bH8cPKm3/876K
IUs9XLp6rCWJAcQs4IkcFwrQGasOZcb5h58RFFS3E7hOy/FlzO+6dkl3K9azaXP6oAEkfcJiiHWj
x6uOWVy6/dI9euESUMJ4gkP5Ko/OOefJeosX+0PI1U2AeW484XiKSfgs5xUwbw5lXLmcFpqM0uPa
XdKNjyw08qXf9AwzLiJ8hWmclWGUpsPikLf8+SmwRBUomJI0mvfYZOTkMjMcJ4ny1ZssT1OCUgx7
At05TA7WTh0GApFk4mVeFXGsqmJM+23SDUoGem1VT4TmeifefM0AQghnRfwxDUFS7RenRTOJUVVg
nm65gEo/LUJvNHMwoH6g3zWKThgNWG5mlOSP4qVoCtWTriN6Y9hY5aTSOPviXru1ExKagzAxQwSP
WTGgtIQlE/8kkV0fMH1aRZyUwFpLMANRteUhC0TeSAIRiH0PmqtorkniBSUnRjxDzP4FplcrL0OT
BUd1hgjO0UTscQkadxivbMP9Zy7Bab4zL4mH6mfg3dG2lBRWRMC1pHUBwarGz899GYvenoT4MhsN
DYKI8rZSJkdsPauXnAD5cG9vb8nGk+0c+eVTi/cbh+LIFvL0CVnYzSbi7GaEajJ3NaTjW1w2AHMG
N08ictKWppjwkfC5V8xnCwvbRQnmG+8nlTrYiBLo8IdIP7qtnPWegxLt0qgUXWZ9fZUxV9Tc6uEW
WMEkxrwTC1ND+lAqIVmngCn14+Zo5xli7aLv/k1JEhbKkl183fLK2ZfiQerlCsU+YPptLSkOqU2M
pZ+/VMlIHLacRaoWSu0vDfnr7PLgVp9P7rDTzPQT0pXr5yI7+xq9bV01F4Qnp43h6HhLMOBefYkZ
SO7cHstwb3CuNsU0LpJbbc3pPAxBLXUWmPQD8okm8ucMueyW2XJRawc7h2yjEWWVd3bZ1L0WrS7G
B5yuSRdNJuF3dI+oqkf7gmW8blfkZEn5dxqc6wEHD85yqgP26DiSDVw0plV74XCvCLCMhNahiVVs
PYQlzKifvR3Ki7w87/d4eBFDQSKJqp3Dh/mHu+O6gpsF0ANhUlm8Q7UJQ8PS0CVcoaK8IQ9tzrrw
OCOpmW5Wz1R5f7KX6WX1B+Z25XtE44nZPPsBGhMX/lvRE5IHmim524bksSVm91Et6GIW8xJddp4Y
JNaLLK8ejGNi4NgTw3hehzY/uR6RKpokPULHBBHjfimTY01TwLfNiMusG8Q8sd7lo1uuszbhffzk
AXEhBGim15XLHm62zOvv9Ag9brDsXPwC7ZF5OdtnRHktaHHsvxODp/9rxj6nHwE6yXwLTv2omaT4
wHQSqdheZyv4+DBd0Y+TSP+3F1HC/VLIt8J/XC5ERYIXKTh9S2znmXBN93QbqhFQVYV71Ku37F//
ftRRr/RKXzYa1JL6Q+kuMGVOTFxjPg7FE+YfXHidFSQTYVliQd76YsANpuComYBpeM7h1C+YmmTH
qWoYUrv9dBaRfYyM/EY6u2X8yiEXHswxOhCKS4Xll01OsJKpNOn62vj2D6Fz+dyuSv7BUf56u68d
PWhdGKcr8LfBExo9A5voMRyVnI9ohxhFtKh8lMFKRC29AxbRebGBBMbRBBbAoULO7BnyxCKuY4cw
kGrg2jjARO1Dkw8Um7dJskLk1Aq07u1C1UTW4giNSr+hBxpQlFG88Jthu8MKS3VsfkqWjMnRtG3q
SRfV7z1ULk0ErWy2LXKf8Vr+A9SZAG+tVZDglHHrFmszU6EXaQpdZeq2BxUFjLH/x1IQU4ipNFrd
sC+4oXu45Dgzo8GrtyrHf2gtxZLEVECxhMsTT6oLcnteJkpnFBffU7gS2ijgWoiZM161ItdGUPmj
aJ7kORVshwRnC9AKPdGOJxDObdQSDJxYCghODpIKolRp3OWKVqNoxCWyaFm9HZfMqjGxD+e6hR6t
rLnlVqMp3PojRESVbpRKYSaseWskXCEjp6LUMvyhIbfMDrc9oY+g98OIsGhpXasgJCwGJoV4NuCV
RIxXvwRz8hDAMwAg52lPkgfvv+AAF4ZLmhNgGvACcWF84t5NLdukoO9YTJY5dlZLK68NNYcYeVaQ
xigCzDsyJhnVxlyCxz2AENdNACifYZYv1KyhJ0GzXKzx254uo96d0NDsRdlYdm3LCt9obkFlOo/y
xrP8rq/4Puu83TfQDXiCE0sLv7L3XgeRfRItJhoNmCfL2IawR6lrcpiPAKqyan7Hlq1JW7E8aqJS
iD/f6RAldZMLw3HkWOBgz4PChyzyTILQfVFDVtpmXVwCpeciPFyeDd4pkyFfiEEuW+8MFhKwnnJp
wMdJSWKY52LmJO9pwbzvlE5fThOrrod0M8+Ta5EkXF9fE976l24bHCYxfiSCrkD4ojtprYD3heK5
yZcY5HjSKKMQK83qPknlhicC2MQcqZPTy8mldJNYqRrOYP5zzRE0O9XQqBc7akDJDKtnchhFSxQW
zLKy7Nodp+SJQOCOnBGfo108k15ijDo1m9QdclCgvo7EZrmHLraGTuUULXRVYOPG6IKzltqZZZwn
VbHj/zGIW8OEMDApzsKoiwgVKx86rHNiNmUnXEuRUgHC9gppR6EXKNyC88jJJPEcbmXERKukZxl1
fmoNotSuQe4yGURoWjggIZUHAL+RCYGTo3/KzMRsUQOnHBKRe6w5iWbNYzemARff9pc+mX8qqfhP
s2KQNaLYz8iZAxCAD6DSRyTBiwV2G5Le/kQv1fVDLCLTx+M6puPBtOqnvHZjSGM1I/xboKN76vVs
zt9FySV68ZUsTV5zU+l/WzVnzxQr2YgvGOYNJJpBB++xCjSFwtT9Z9iiOKQEMP6oRi0X8ETTmuNU
p0Poq5aIqIXxIyJeiUgMBR0s6KAavMJVLqd2lbblm5L40Lpq/996ysyYjeQJKsSDKgONEJLC4D4a
e30SXZuvEe5Wb3pOgSCvShahJjHlFdrI9jff4jGsdSVn9YDClOhOcCMEGe38upEYML18Z6BWKyKk
mIxLQLNUlICHpcFCEgyHrxwyJ/aSHLY3EWnk2n1TmhPtQWsNnVHMKfPbF+WcVBqRNWSPB6Akv/LN
JIyJpPGC8DMD5eUOKsdGeclt2V2pUoYYd8RkC205Ut+B69/n54O76bwfcEgWJF3IyN0XOxIUJSV3
7FRtWGJrcp7/mvJNnRPYExWoV/qbYf0nxg00QYWV6iqlvGwb9+I0hfZHtUK34J0Y/IRSBHzo3GXe
kTiNhZ6wri8HpEXbkuzzLYiQOlb/xfxItnqFOwpNq1UhcBbuF2gnm/8Ef1p1cqGLNJE9T6j67t+3
SmJhck7doPeCl4CqiiJM6UA5wqZpN/QxmGNYUf+r36yr0iVTUjeaDEsVpev1PGbW81KS6+DrOfN0
gmYCxqslYUkCPnoRdvGFQaK6zGZouOsWp7N6jc4XYBpuB7Dpk2SkND6YJXj6F/+CnyGMcS7LGUxT
M0V+46b8BYUOY66HIlBOcPIhn/+xdfqJ9QjyrJKq0lfGy0Dcx6jM3iOLLjtu0HOVV5MkAVuj37nZ
BzKJS97CkFwaFYSpMgGu7YS+Y/6uQFBT/t1SuLR7t+Ikke6ngja6kb0+NTLnmA5URMfd2g6IbVJm
COmJ4q579hODlJb0owOXGNyfNajnSZmxxht8hiN4EbFG4ue3pQw6uPc8izmKxzx7Ch5ugOvqy2NP
mRBF9cgqAtTO/Bp9BmZbrEk3HFAveouCwPs/AOJYPSXDJWP8Nww9QjYMTxuZg/f072VkZajHWJx1
8ExJ/KZiTSqex8aN9fsf1PK4A47vqp77jMUxJsQSKzgtfoXT9XYXybsSgZKu0G8XqljU8x8tj2CE
CHLCVX6wIayZm9cLZKdr6jZD84KENLsIpfAXfbrsa3L2Lp0t0iSfW71dZ6KJ2DlgJxgGPYFmkyGX
qgFpFFXU4AlkzjFvz5FRTs6bVX68HpoLyY6tZLE2k0GiO9Fp/WiSpwtPDMEd3PnIpzzusxc2FA9G
lqfw7EIq9S4A9jbJWtGy0iPOWfmLaNB/Gd51LbU7UVlnLZJaCiyBJWiClOE5DLBC6TWf0pngv1Yy
Kz4/ue6aZkXBfEdyySCH3W1e6Vog7ESpySCiec8X8UzP95/GNTtxBvuj4sEkXQhcsjTl3iRV24Ce
KjdZ2D7jjkx/mOsnhxdJXmMOSJyY3y/86XanB06CbW15dYeQMFp1TAWBvLuLNpZQpZSFPdQkvagi
wfP7AF9RBAtq5nUAUIdvTCmEk4RVyMIPoK+j65nITs3VQRi6ToFr26Vq/1AEUcl1qbDc/05mX7d2
G3ahzTmzr+eujJPnJJBLgCEiSl0vz/fIqUOClokSt+uVChaFeWCemdMjJN5r1ruauklOIjC3ehud
J+ed/+oParChBj/ZL+wZwWl1dZ00YkCxA+rqa+/8IiepTOtE+6aorRcwQ4gaxjq+BhhIUtR9iOH7
yI99w/CQz9PzOGYdRtmgIH7E285lrNic8JrJgHzl7HSDEZaujF/izCR7WzZQnojpUYaFnNc55iA9
o0ODD+hB1RGn0qxyds3oG7OMOZdzi7/PNZTwqYYqOYpdCqRt4jPe0YxukjlWrT6aS7qBndhssns9
7zBnnMXqumckvZ+Lg0N7Vq7VG7POqe2eN44pu+1euYXb0lhfMyfeFOlSMbrgiRWLPKZsY+AkONgj
5Bu0+B27XZqzrXGhPxvzYMPKt91p/nHKtN2KqweuJVKbt+Ivlsavz4QMGeU5zLYcqEM4yGGaWR0d
QvnpI7FamDYabxYXDwuGycXvZpILhUojZ5nj3Zz1cJKx/8wEdtXKWlRDEpkixWdQitt5Imx5pwQb
W0gskkfyYtyf3MVcwS2hHQ9NueEgG/yGDGQt0ZNUna0KapJYIcIXOpiKXOJA7d3YEUH2u9uRUA3V
rYMRknFLMP4uBnFpOIauGQDk8gOemKjiD6+1qt18isbCH0RJEYielezHcO/MUPgI+FTVmoVgQYU+
koFEjyFq8v24Xs1ffz8P/k5JKIqb6QUj25AfhnxSlOtDx5KZ9A/QDAjP7BTrBanlXLZNdCgxLcoA
hHJg4eMOHhcZ8IMRnsDx0IWSnamPnyJqhD2OrBfoEAYQbI5TorSKBpYQcEoGmfj2AbGCwcLqGieP
3wp3FIs3EYU4S1dlqoyaAtu0oA611qaZKfAAtd4wKC+iQwo85IOulrOavAimbaO7zeaA8/n2DFzx
bQ26cG+teWhqt4Bvp7//5cW10EOij3vUk9g/lmnpaOfZi68WTU1BL9gmbd5Gljbm7eaaQeDYgOW2
SvDpotEnENYaviUiacSPaHrBRr0FRlWrngV7YTcRPvzZeEmPS5L+3IOAm3vsHwqH2RM2B3qMie1y
U8MaX7snixdKV0/iDPQcXkSfw6iReHpiL2n62LrEEG0LjFQ7vxeNHj7XR1KGw+Rq1wNFI78cM0qg
D+wXQbuzKqDuyN8ncaOEwQPqDZ1/u9jtJ6D+J3cc52MvAo9dSoVjkkNiZ3pxvozkdHRTACNFZQXY
1xOtE37ZXlbm+ogvpJx9SdgAfZdazq0zGDtMAwi1vplSr9v3LoQUmZlKs/acJUdEuinS/LctEZOJ
oh3na/h9FBBQyAwifPhCPyavQlHqKopiT3clHkc+15S4vc0TfDZBLMuWGvfXcH7v4PzDO6ImPtvy
N1zaMpp5DVRZEJDe4Xd3xfD84rGJ9r1io3OTzOxDjhHw0QCxmrp7PLM1FCUv7T1e0IrA6wEZH8yD
nNOHdsx8iiwWSI3q099+ornJX35csva6snBDt5YGuuuc9qVgwuf4xYXhzjaGwww3z1Pa7IbVbUTp
In7D94QG3GZfSZAnY8vx+8Yt575vs6BEdNdBN/Qxvv56X0RcUhkqi48laoxdj11LPAUFeQElNhcm
GWkbPH+l19l6h5RF1OKebnePBSVlX7mTSAMS+kXN8AMst4kDlRGzES6sS74cPZFnL1cPc40kQjAz
hlrTwPJgvsnGTSBaP0zOT/BqHEYaleLelh3stkH6LDsUCDdViJ93YUvRQ66hwADfaPfkMbamP5VO
x+XApjLwYZj4SiW9TLJTHcwbiJVI1oVahEtp3BnV7HUkbPY622FJvUZdhr07z8UphTklsJUK7abO
IPanhjN0QVPYE2FPFEAac+xiUqY49bEtq4tzZL3hzfzd9Z8o1mjyIBuCx6RGx9b3xW8ofv7AJrJI
uO1hH9ML9V3kolbwA7eERSWWFpq6m89QZFJ7CJMU/6/SAxsLo+OawLlBHZxbSjYaHv2ctZC6LHGU
kN684LOTxhjLwTr8C66CTtN1pdLurMDvWn038E3XS/J1UE812fTw7DrnHPOK3D/im1NAO9efDBGS
K6AqDmZ58YQB1P3SfVXaq/Jvmz9yVT55U/ndqHziiy5xK/fp6MF06jlL7vGHK5tV0ccT3KmasQbk
fTgb/9fsKJ+GDI/lJN66PFzZj1QVAigMXAeWoU7861c/sbjyUjlt/a1nFH6WrJDtmPy8I9us3UCg
dFtxb+EDPn4HlmVxFMt9zPj1mhBJlWNPntb7RDFpKpbHDtY6Nh52LloXGZWLukpqmigWp4903JUo
i8E/6dr5oZa7opnkniaw5snN9jU07v2DfLMJBJA9GGO7SSG4J/w+Xt4lz/W3gNMU7S8aiLFAm9XE
z7tkBFSLAFlm+w2rb4D3t8z4C8yznTyJnZ7mMZq7imxkWxSvh1IVhVyJy+TLI/NMWHsdOJ3d4QAv
abSoMrGgnz7rYsMGOox/4U00X3Is9lDkBy/vLA6PQhkPW6m+S40PThLYyeHIlPGD8x1v7t92T1I4
wjj2DfHU2IPK35flamjRNT8AXrSjsMC2jtCZVB8I7X+Ul5BHd/wUaypVXFCmQTiCsmdkfa56a3/X
2xfvpqYlBLACUYwKD1BNdItvyA/25pSrNuuPlUoE//V1tyfi5TwMxfD2w6InkQisPNu2KYjAKnlg
9f2LCyMnJCDqtikXMnHhCpj4YhYF+1qwf3Ne0lloH/izwhDG9O3Gp0ASdOl7LbtYyUlXoBmxuIkf
TEsG5M1nrE6S0Yh1LVeE0yRW/rGBWpHtSsaAR4vBl1vu00w6BRu7O5JKJXwyGUTGnjQQnAFfpbB4
A6o4StzlwKn0bvI98EOssKyLPX5B7uD62Dqv5rcPcEorO6CctKNReHrHcyueYf28Ow4becEMHrVu
nyAb9iDnSPjJ69ogdz9abRjSyUvi/JSUiCUKeJaEwH6myvELzoNhvvV3Eti/Hc4no4CMGZoot3En
WpMlAI+Cp4xy2eABkrzxCqUzrKdExPiPNtlUcE/65yO2H9+Qxb4RwP4R/4f1g7lQo9lQh/tbCTSt
+YZRWDAxzFu3FGGSYUU5S5KddfC5JrIRQU4xZO0QgZ9XIbDA0B33yZKIkPwq0e73bupiO5VQX2J4
GKiGWaYcC8yWzxD0YIZUPL505za8bzULbN3nvguv1PJ+XTa0cyP4/NQzcqxxzS6TX5tKPG6dlzRS
q9CLFbgg6AdspzZFWimwI+hXZ3H1GAor5HophmNa0fnjand1uxo//KBwBSE1dz9VIYpc7E/I++5K
LLjRCTuiHzJj/XLaJzPGEnr28FZE1C8XhD8AhsbAgU6sG+Dh9Vl4gdnJllIDpEzbz+vStCb/8Kyi
6fcA7p2NcrlLTUcXE51jUfXuE8EXv/iLA4I93K0xWYAPt9U1iUk1yN8emiK95yml1f6S/hBlOCII
MmvH4G7cslDDJ+czHK2vEhHVzFfCNZm5MSABZpT5O7JY4rzoEhOlG2ilLnjulYJdAYWdG8l921Ew
Cyn9Ey12tvSzDm/5Q3ACOSDXL9mcLUirQ1p6QIx1ZRTVq891lKxiZVyYvaJUN7HK1eQux8DGpfYC
JYL1Ne+8DSdtDTSiwaJBKtRIf+xBh3bTjeozLu0dsMa9UE6bNEaT3DnX0uacZApMlozI/hh2FDmf
em5s3g0RleoMd5YrHb2xjptVcxsGANqC35HosM8NY7BO4ro7fpgFF16SH23oUm7DG2aLX4XxoB8F
2hfB9oUiMASLobTj/twc2Ldo3UE19tRGDYOIfwoyiLMd1Qz3Llf43uGjpCfAC2uGErhPUQTUBggn
/Tmju0vVbt5rodLUIHiazVZ69tNOWZpm7aSc/TXglDN+wFlrrWJv6CPSsdp3vUXxQxL+pVIw01/3
FMVaPH5g0O3nfdrkcN873qsGQCLVlNPfXVr0gigxKTIY2WUBFJSS3Bx1M9m7iPxdnrekCrZvBBXJ
ejwEI+0pxNku+DBcQhWj++O6XhoO1Ve/dekxWAzaWifcGsCWSTQOzgk+MV7HZDdG7vWrtI7PqWfz
Jg2y5Vzy+3DbUlHNinqFtY8rFcZGUBcZq5MFIz0xfsrXgWyJzyErk1PZdPSls/914zjuSwOC4r3N
ydvB7KQbb0tNxI5sFQ/3Y1UELWjtOLtoIUS9sDLvXQqOxQTi/iXcP6rmtqJ1zbq/n88DMt8OmYhW
A+7vzBoK6QXpH585mCkuDd08LJJjerTLWCK7T56dzQMo5PyBYP3vIsFYftD8HD389yZw5DbbtyWV
o0CPr7enCGmx6O3ubqImqRJxEkGDFmYRyJzc6zbub86/9DNAxqRIhiraZ+Px9S2v4H454uPCLxOi
593s3KXCJXWw5oUDyQ/xygYK/Pb6H2KRPYMyFeEOiBAZmw1aRG0z8YPYh9lpvZkm7zDKNweNIkSE
nAyNn/tPfEQid3fjjpL1gaZrdH1cEPiaZtbGCmBHgG4hvN0c5pGOMDBP2zBL870b+sHr3lfzelOA
qunKpoFciKGllHCPo2GB/0L08XhgsRkwLhur6ykvshaUVl64DCpsZy2xr0wfXAWyeHjHhRc+n1Rv
MM5hh6Kgszd+TcRvOm5GWPpTMp5RJfEbDv49ImLcgCYFGCJg0cJCN024yRZHRLi54j35vM8A3ant
bfiY+8MyiQ/DTpKTUo5kPCtCqQFuxNeltsbPX/AATaG+0mE6h5Xx+AMesi9SryYP854xX7kaRNx6
GqFE4U8KVksZmwYUw6/tH7GIrBvq6Ak4u19bsd8y4gmjTgONPeAWB4QF6HNsEgK8zcRI2CZpAGhc
rdLfI6xSN6h0W79tMdYO4mN9SwKQx9u4z4UmJOAr3BS08qxYH5qNojKiqHi+Bx4vs+xteEHe+9Id
bzyjJr7q7JwD18j7jxH5UVx7PVTizQcslx620oXqp3toyzjG80AQbrTgViObxzm6fAu9XDcoswTD
sIvQY5swD8idx7bEmHZqOytyvT7jfu5lzy5YbHZDRAGCt03CzyjDgWy3oLRVoXyDwn1fSz53/XGl
AbAkQV8tfBumzPGVady8+tpqxIYkjEXX4YDtOvLp0J2FW4OOZGJyLlSGWZ30Kr3IuS97QXdqYs79
Wps7xENsYAlw3kttmrqdyHuC7lNqarfl6xFCYTIoZHXO3h6Y0J+ucVU6evB9YQ65+e6B/CWa0Hvb
5e4ClaDFeHx20L6DfjydPWRxF0ncMxlQvxJ1jASe65LfZTAi4fPzNWcTgrfSJFzDWIMYBN6VUXzZ
9obK97+tmjrCw66SSV/npj4Tqjk3e+IdeWH6mTxUtq6yOKOz60KYFAyUchZJBd6+EH0xAnr6iTbr
fmQZTCxCDxujmioZLg1TrWz3CEcNremQQOoTgBwjXPvdqxOfHoEIMAh0qTJIM5POzL3CIJuPQ92E
jkiBNDtNpqRYxPasbW177HQMZ1lMqrk7jtPO0ySPwUQrYFhcwCpFB4501D93Ny8yhx/zjK3NEno/
fSIxFbKVkQ94rlGUumJLX8OTZBuctAOmhefRLNTYUZxNlu6EVg1fJqOBPM/jpt6ck8k5Nige9IvW
9EF5bp7PG1pKld4L5s8575AzOIE3HA49cBHiJY0aNPmMbhSsS1Ld/p6umBe2uVbB6uGFqJ/ijVi6
amxS4sbevSA+SLpJIbEn0c8xQ5nQBbesE1MIp85qTQdkBcDxcisJw2edlvolojev1Drzm2NeJsNc
6e5enaa6YUVAE3+K6PfmqxZpRZbHGkdoi06933hvmgEkYaD9t/zShzREx8FI+3VhoyLGK1LaBCV7
Z1Fx4HRMUf3xvoho/Ppfgb5+T6sRj6ynq//nbHzI897/PClHNnoS6Bm4nuJ0+VodTUeMjXaYvKSd
z3W2mSfTthAvzwfQzv2h6xpznlEiB67QuQ6xVauunBM8XF/NOM4VMvKysvVg79x1gwnA2SP4KxoG
cWm9h1rO5+cLKVAxNm86j060IOPnpTUE0HaAqNohxHio8NgHLkOzv8mAaGfRJQypUrg9d6VLIl6H
3+1MUZzpCJ/BzdDWtSOT2b3ZCpSq8TRsb9dUoVlJBJFvZJSBQjt0rMK3jvSPOskrOHEtjD8qbnTL
DuybYnj5fs5JtZh/Sm4paAkpqQYZIdBERhc9zlni9eE3Mnz0hXqhOOJxbgo8/+WHXyKeD/EYNSTT
7s+inQZUF0z1gGE3FAAWqc9iqjvZdNm2n2zxbc1AejAKL2lu0D47w2DBSFRpEnnsYfLzxEbF++Si
+72MlFvD3J8wvcAjPtHXk65P/uEuKLumKN2Bg0xz+dCutTYpGmAYGQYFigusUad5zyUlyAmgR86J
HCJVl8iwUjegC0JEbtXWYjze0D1Xtez+SJRMfOHbM7u3lBBr8tlxwMaqx6NgDOANmjjHjPaNSS8Q
xXvE2FPaPpHAO9vKgHvRPTnC6+ojCEFzxAj2/Fa3/C8sO9w3Z/Z4WtQOy2GmaeRFqtlw9hBbcyV0
MJUWB2LAGEIiOooj4qBv3ssovKqZ/Bwz2vgllyEj9LAId2eBvjkpaEXwiaCo2KZZOy9kic6+zqmD
anodo+e842X1vZdxMP0ITJU59x3JN5s0Pq1ecMAgg7wk8e2BMH9sj8hW0NZYuajmAILBq848SHNK
vKx/CSxavdUSCqkbydFce9+qaw3pNx+tMwWHM0stn54mIh72GJMp9/IRKc+i6JVjjMFV0FZEyA7Q
1brelc5bbv4PgsS/+pv27tFxCw+zN3DcIxo+s/6RjJz1kh7KOp0w2EJQ4zbSGRUC+9P0RdnrWVdo
AQLX3aRCsXZ6Cbj2Rvy3zjoRK1cLdFq4eGDaNXl5O/MKT1zGKsJXPDJJTrfg6QPEG3ExfmalgPb9
ku0vFhhuXjozOiRvK7v+nLqw5sZuMBi2gBl++7aN43FxmKhJGbTpDzzb9TTjsO2HB38s42SL3f2w
DulEDZ//18V5CbwyjIFs4esT92wMqtckCKWLdwoYKXbWtAIe4wxGq1LncHXJBE8x3Z6LSB5vfPBn
mD/EXeQGZTkuCXHSkZX+6Qpb0H4h6E6Pu5AZifKqWN3pWIF8vPm943lSk6w6AfKWSRGCg1+ZiDVu
n/wJaCRK8cZMKWgP3wJZuTTxN+T1f/Te5bs1cZpg84qtCyLiQfZtfzDcAztcg3Uw/T35QTn1icVa
C6EIMon7iEnB5y8G1/DFOO6vCmW0CkaKj5FtalIY/ia8kv9ai15dR2RwDIbYviSwKR5K+wgitPqJ
fWZJHmo7gMT7GMZyeJZHcMV2fAdzKZ4rHHvgRxKJCrXysHx0o8AVqEWL1Nakv4ta+/T0IMH0QMMi
nLdw8L0FlJhCDsbgfAIVnpIU8My0fK18kEciBxlW2hkvWk17NcFUhgqkd3dXStFmqy9w1SjHiqTb
lPCxoKVv/JBwe9hbGZGxoikKpFTSW+QIvmiiJT6VUJFglyK+s4au+a77xdKQI/xS933N7g4jBtq8
mvnXurjRpQT2iLj/XpoYt+EiP+wfuf5/bpkVLnGG3S9I53dvRLXcA/3wCx6NkgbMrDl/qynvzxF6
IbA9bYCo70Xl3TRmB5fKe74/+CAcfYskm86M6Dilh1mR6g52clISS35Hnk8U4V5lNFH0+etJFO3Y
r1mZjCGku+xoclR6mWysH1TDpdebe4FEBfvWbWE6KJaNkbFg43ZY3iDQTtKPxaymbnwdHbFuvbgQ
2EMo0mzCfi/cYDvq6t09u0EOcTZexqFxGpog0DmpZckm7BApMAIRhoZcsh8fn4/gTmqW8QdRWptb
VWIRIisb0W15kpd58fxPi8nWEuomnBY3ubsoDUGKVBVM4ruR5Aapz3hEL88FcDhZbPNirudohT4z
E+uvYaYHTRRmaZuiXqbLxjdtJNZPAE7v1knnzkFx2u6VEeeDh4tfYJDHls+0ZDnFt1x4/n+QR20z
5tGArKonr8qivzowMepZEuNZmOlAQyUhqxn3BWOmvsxjEfkL5B17y8ceZ5jGO9dLyOyDLTvnZpz8
c52vb9F9ndB5B1g/KUhLZqt9BdMU0lTpHCGos9cKyJZkDieXTFv5T1j3Vyrs9eozFgkpNvDO7GWl
lDM19lTkG7ZBTVTQNKkVQkOkikP9GvpNEPTF29cPUtmVdqkQagw43wLtz1CyyD7wBv7bPgAKq5Wz
PUFhLHSR42+GGRzcKyCsy+7AJ6INvvA696E46k0CXnW9BuxY0kjxIty6O32hoDiyRDOSa3Yr9pPO
PNvQOqo6tSr4PPrnWaONB7pwiW5g/6UOFL5xT/BtG3ig4x1XqnhZ9QYi1VsOXI1dlT73moFgce3w
dQznd3xbfJgd7nv3i1cYnpTCMdKBlQvSeABodSXsG8I+qX0omFXydcAo6+e3sBtJeNgmW42j0jxj
ovSq5qvhnz3SqxLUpnGGE4WoKbi+U0lvsf1uKtQADLqtOnKfMaXYsxVMNTkyZkT/J4WkESGE3Kth
CtV2vP+dzlhKEHZH6OBGcbEDNknZCNWuy+yoDSy130mMharh5k8Dj2eV0i2RyOc8eoRYcAFzwctX
PerrX4zyIwtW1mOCJumAUD5qEk/FbVEfKpWjpCrV6vO8q5z7z7PdLn6Zrrb4oxwbWM41t19yvnhb
tWyo34PyPVLm59Anr7kTH3Ul6bkH9qzP/l/1XZtJ8xnyXHIgXakANNHBv32qhk/ymutYIO3fdL5m
6bTIp4nPW4ZqL+H4kjDq6hViRPCWHGNHKY3AnOKpesYEOHGP2my9zkgyib3nDA6lgFbefvEZv9sW
9CbV7F02QIGXAAAnQ8PHmP6JF0c3IIVxZ5V7vGDbtapI4a+uUYlmNBGndj3t7FBbW6JhfRrIhOg6
Z4aG4iGrRgSeDIkrHBFmcBytUb19CsbDEFVmobYL9jNjRtCg20adLEEDJnk89W4peXKlBq5dEH8E
CVJWpb/wG1a+gCui7YxxkMfR3d7GTAQCyY1FvM5ySYmeweQBgtTxNUbD6nr0nzNBVL8cMQmIqzvX
dHugEzLvK8u9mm6IPoVIwSwkgBrpuSnX2IUfqrdqUBMqu7sn2unKXbWRw3C4enh/Gqz0BKY8Taai
yEoYX2cYQOugmN0PqyhaOlwok9wjo9Tjj70E9o3lKXIqkUcCLSUVkyVI9ZFWaCRLNd4gGP7Pt9yT
6abgGGO9JlrdFTAYETuD/6vl1t0d+gHnxSd+XjRKRIO/PR08j+kVMq9vyEEGE1JLtu0BSzITvQkO
E5nXd/U+JfizZYcFRpaxrM6my1ASo3wXrc8zm/U4YNT51Zg/p4pKCERKdnvvKsBo7Tv0fEwlAWdN
oRjWFoq8xfm1GnVfA2noNa1ruiB2K1rLibF1Py7LXnL2GSQtXTHSH3O0xiQ5kg1kMFEHDhZAUWYH
P4EwiBsGLzzQzJy2aKENhnLl2zaaGar2qzreTsj1epVu4uwxKiAcxoQ64/QXc3vdwUlGtlwfszIu
WDqcOVM3qZHRcowi/jVg/vezdg9xszYHYf/UYu/uwQs+E6wg0z/XqXtmH0U/flW6tEOsaQHJ8Yp+
/EMwqKPIRjFCUAhIj2NjB4A8aGiHFIlgZVYQj450S+iwLd2anMIyfssHPpZXHBJjvPDoDhqri+XY
N/x/GjNZk1Sz9BymuD8I+WBpzlPtrU3CK5DA8xK68VnGHMhpq3A0pXWiOyza1ZGFOktwfY7D/lv2
KUwaUHVi3rqBNZxjpuTqBD7KMUPJTgq/ffYD3lbVny7Do259Oxh6q5D7ezOt+fJxRj5gv/8tyS5h
V2CpGdgek89hUxRAs3RkglyQ0ma9ret64dhVBhaaJq8ER71eLriHdhdzBRiKHKKCx4TIPh4eENlG
FQtyFtRQjLjpX/psCOgeINmSe3texnz+VJjtDDgHFPAYitBz4VJDy+6UAzMZxypm/e79e1m0w417
1DtqkmEqD6L5MI68XpVnKjacx08KzPF2gKQByzaWdecMx09HQN2Su2DGQHDF6WvuffcpCK9q7nq1
NmYL6uwDExoRXP4e8T0hDWSlC5PBEHTlm8bol8eodcpHkEePVuI0BVfrlNGP7ZcyWNzzig2E4K9Q
CoSiQmhS7GFArLeXoW8YD4jbdSughD25S6hHO3VXU7ESRSz9JQbGXCP1TBNJ/nMYQ8C6Gci+3uiF
KIyBksccG0kXJDCKlNZu069EcscxscwPTJn+T/4ZBVamNjR1gdY5zdEc8m9pOzDyINf73dHoWVqn
ckGK9Z326MRFjDdOcZrVmHPPvnYUxfJbPU9yI9b5Vy9knr42M0+I+XvUF2AOMbJe/uK1ziK4ZY3Y
TVEz2CYV5Ywk4wzc4nPfJbVChoMgyNpzz809r5n8cmZJ2zif/Ss/WhZeVolMOtTR5SoHAXEyXzou
Oc1v2kcc2yUsyOpuTWT8LPFhBc05RLSrggIEFZYzXCquLTwhispbtEqUDzW/uOz52L83YvAXeVl7
ixob72GVxHf8LtQ0sYR+lxJwuF98yRwx4eLAWkGX7ZQ5Dmmhi50hL7Q6ecoTCPAPtO8F5mU1qfC9
ZWPKeCcwE+mxgAj2gMt2WOlz3JpLTAb0rsKnJ5+nMx3Q+KN+kMyqnyi/BN8LgQrPMcO1kF/K/WRf
aMsQT9cutPG/Ge1eG9xjjuZgOvoZK19FdVyOUa0cD15CmE9TqGyS67Zxx4tLS5owTmKzESpY2V0l
zrl4ltqNmd3D+3qjXDlnwQP3+kkFITeIyQIsrk7V5dur+xQT5V3RNgRaBH9cgbvqvGbCjKUP531q
Wp6JDOECPLkmp9jdcrCfZ3tbTEClYisKy5HfcZCMrJJmo0D/H1Cll9UQgD+5Ke7UsV8Mf/HVum7u
lIMkcKIFcyM7yO+wcPXwu+tM3s/99IFAvXk3XbmSYywTEJe7hKlpVYSW8f7RxLaMd0UEDm1aYwIx
R1JT5DutmUG6iWjvLRp4w9uJeRVYEengFGZQPHWfvzblobFFj51sWojCetNxbWvco6KlVXNpr2xW
wcKv8YZbsJjqtIB1ZfoXC77TkAjYcv6OFv9b7RezbF5lU04t2JEGAYd65TY2vqfOMTaFelwfV/F1
pf2GvVPNkpLc1nZn5pLlnB8iJ2A219eCZonDGzlRtxdSO4XUQBErLZHEy6mSvAN9+lW6qWU4vEVY
xx4/Pi/Ahhb+tCC/fARDnhsGPP/xc6+epb+EQNPwgPBD39xK8WOCQuBnTEP92dPvrpMl1HPKXlF3
BCTmmyOJM9nHW8MirKOgfelV/SOLhr+nC/uZaTRNAYIztwtMAkk9ps2YunHq19GMsqKQoJtv+VtQ
DFKxHt23DCMPwq96TJ3VaM1VlSwye3y5Bg651Oxk0HUW7srkLbciDdfKm0iuZyKK6TT2QbxwdPRb
Qk02WpOg6+ue1gJDYTu/5BO0RlYroPO/PZ6LTVF73Xsy4ZGygUMQbcJNSpqbihVpFuwJHsAWVqrZ
7VM8+Z040/pJxxUo2gs//TigoDlNmX1jruG/c9e6Wk4WI9JJ01mLj3FlHZnxYW1SxL+lMnqPvUHy
pGjOgOqSSBomEfVX54jR5dz6WsAbMxObF+9ls+0J+m0Vz3RiOn1WblUZxxLxA8fhFZuHNyYQ4a0M
PRaUY9SpN25MzeTxwjccZam6+36Mq63u++TH6iJEUZD8D4b69P04bKTgbRHDNWA1qD7T1Aff0jA/
RrgxYBRXw4IL58/BB9Xi6N/9n7V06i3/iJmldLJoIsvk7LiPqWi2PNW7tR5IJnzbsXK92/3ckTyZ
9vrBoLx6G4MU7KO0jcBreZ8lo8aQ4zJ4cqjTmOABV0LBYQ7ryViedo0p3/Ng020GCGn9Q+BSdxG6
pomlzaxC/7z2UJx9QGPpjKYaPWfYQk1USj9bH7HtcEfi1MwGRgLCRey42dhhCnJmA/wgAIfo4nSB
CXV1iZMOB20g45jaTgZz46gq5+2AmcMLXrKK3xlsLbde2WlZorx3rRKg3QCy7YwXL9eYkStWowLO
cpn7PCpKdd1+PFLxH+KOG8FRIvQlKFBQ0PmXyaKxwZE0GXUxAKBl+cPc5xNTIkFBMpraiP+OCFnG
1BPnpqp2KHk6VBrB3lGt5WhdjiKk6sUYDQ7+DgQCOndyep7U+i9hERY3da3zRe1z8vadRqM8ALrd
4Kys5v76RFsrr5tWt1fLPQUsxR78UzkfhxBjCfFOFwm1yH87ZEzYi6CJRMll12scFwmOfJ2W+jDu
yk1am2ufIz04J2+9sO0F2D4ICjA4lYnVC9GVwm3qrPbwp4k9IUt0SYAI42kAT1ebCbg08pb/A9f7
wR4TyLrPaYHRW8NMcJiChr09W1msQJEEq7tZFzQDeEOKqyGFABUaOGglT+KDlG2E5oD6QQ+PbnXV
v0IasABtWi+WNHESPmaFV0EwFz8SKfnRag95Wyz8NckbXQ+NiT3i6hgHi1+NoIKWF45pSOA2RwVv
7A4WRZfCVyI407E0q540iyh+yI94+rWT2EEryiEomUxb9GBrihG+WjkdJtC+1JxJeJWUj8LGkqQC
Y0AOjHjs2vc3gv0uHmieq6aUeS+WrpXNFh2esyGWse+6nuK6McHxVs3dvZKSI/VGOQmBpJia1/fr
NcSrsvZmDO6JFOdMnVzBDks120HAEpq6vulqWOCyXWcT6BWUcDp+y9LJMMfzy7p1ND94K0lke4V8
PiCefI0ZlDHgmVtj5LAI3Drlq2FcQYG889XARfeKY45wHVQKrgECHpGLotUCUNPMqGhhQnEavYDR
ri7M6B02CGS9ilC2UeXTzWl0BNm7GP4JkzuluVX3AiqCZDDXRtZwbCnSyAMG9jBmCvctJ6M479tY
INYemRjxQmzdBiUu9lhtxlM8Zru/AdOGHA3k+6A9cdiVBzk/6rC9TIwD6u3FTBR2YTpNwIAmRS78
OHsSb4I96+RlMNw1xShmUF3DKCYX/7FyyKZMOaQHnWB8IuZBrqqdY0U2t0WiLg5u4BupD2ZxfBxP
xZdH/bss+BPr1adQN77tDl0C3AlRvwOVqTStjHRB9OK0WSkq/i3WX6236vF2DuxbDwQiSnNjWXt7
xQ/g24LEl0/VXAQVGeN4O5d+Foz3Qcu4+BenLn0rYKb1mqkH7sMuVgrvRaz1B1k/YdhH1PMGmOYx
y2BLdH6YJBse3O4knE2uY8H3bpKJt+dlIdL8+IlR22Ddosdy497imH/+ZZzXu2uir/vKkTJLbQOG
ZeibwUBtmlClWRJxTC7G4S3/hani+WTY5FXs+bPCn9iK52rFde8BDdFCKww7xBL340ifj7nyXCm0
QXbUy7s9aBE7+KIaZ88VKDobP383A3RzgJhIz73VgU4wPJnZk57yqG6GZq3lm6hDd8rIoR3ds9sg
V21ho1LYkoyT7akj51cauk/tS9c5ka5IS5YPC/e4hHHJYPpagrO2MBxF1Gef7oMm0yP7oTC3EKf6
ljVqh3a7yOfBYjm0jp8FgTznhUnW2GoobfdweWSJKC+WLXEC5yRRgpj6sy+gzNiE/GAO34dnWcQa
Z7hoCjoWga9FcNS/hOqaphdb/J6fGRUJ/Q9NohRs8vGwBJrzeMqAp0e/I9Y6fTyBoTxlJH9bHRCv
q6yEx4b3XO6Fhol3EDRGhsBMeGsu975gHZNQl8S3/vfjR/xYlk76Iv/Fs0R11ntI9HFfFqrh/Euc
WB0U4bgRKNghlLp1TMWegW405WJkq6GCFICs5qiyaJ9WMHk2cI9RuBCXfCn6nNbK66iL8Mu7+kGP
LXI11lwXZZHMWXMt34IcEMS845xUJJVmyfo/jOn8f+KXjLOZutAQ6CQsmS5srPqlj/mQNHzEdhyB
Qe/rKgd4WPFNx9IfD78cx0dHjw3hfpnuOCVMa0tZkMyaJ/jNQvrYdjTqOFJ169F+s4suukYq9zgr
6Xv1zZCspt9UsVOH90cBqABXHCp2t080eYNihH1f2eeHvsXRHhiIA3mRnO0rCuMRyExMrXKPSF9Y
ZfMjehdvMnesm1SbtY60ojmHu08Xh09gONqB41q9SkQBbPXU9pv8wUEu7euVJ5h732TYrGHgMEYg
+bLXQSgye0UzDAaZz0dzdn+gacdHV28V6ia9GyfaNst939KLlSNBQG81PXFPPk2Xd5PiUSzrX0Pt
2oo9/YSxFTpep6vbY1oo34/0xyodB3VoPEqy3Pa/3wXSRrq0cE2gWBDbJexTQRS4AxFMP6+BaM9C
HLHaKABS2V7TmSOG3mfT2tAXZJSqDaJXoPG+r87YOdcxmZ5kbyqBGx6da6glzcQzzxLXZbvkoO4U
p+MJg6z52c5HX02vV6bH9z3SwasuEPQG2kn652K9zBwfNShkAIov41mWRoTKC7xihP18iw+26F0M
3YJJCiBv5UpwB4ZSKEMgQ1hpNx1D8ZcMyOiEybLz+aQ6fSHKZM844wSnt2+VuqCeGFipqZngLOGM
KsJ58c5xJITzrFjgGpckKecjN1bf5f3G4PkM1RZ8cmMfqBEq+xA42+McWGF1zr2ua6ancx1Y/D6o
h8Z73vRXBFXhVg30hKtTAU2Jh5sp/UBLRXDBf56Nys4pFgxtBaAmLPFhUqDtw21vZVOUA2LQoBO4
rjz+dQCXhHHAn8exswuGSS5BDcwKyXcvXjjcJYTpwsyrUF6Wy7HFNPBfQ4e6aTq8Btahul/stjbg
pZzunmfmJQw970RJs55DB4W95CR/lJ6eA1KDX5Uc/JbO3+3yAd3AbG9AzxC0b1gqBJjF3Pt9/sIk
78iEjSPczBKb84v3jrBgwYgMVZL9Ad/iDpQLDix/xd/57f1d8uzX8D19Lddkn8qECvP250FHmX8S
TvPuNxaPeMvD2EG3kGYOkeebz9bvvD3ee9G7A2MwFRxQPeJ26wgWFqjDSZlYQ9nekH4Ng3WYPFqc
YseE0ERCKWqTRksEenVddcM0i+0nzR1937L329/r2XxMhvFo2ooSVSNeH7/R9iPMQ8wnp0dAewTj
UozGsvGeRry+xK85IUeJ43ew1zOBEaK9lDs+IzqahlKzQ6pJlqX67rDtCdIQSCabpwUKJ0nm/d9p
n28E7P5bgnz/aBhDAazm4AMBhh6uL+prgK1ANhYVeIplBiWQS+PRajNWsDVToHgNiSrCclMmSNG0
zDN5KPpHmlzUqNxi7YOty90eNVO5EMoujM86f/HdRz//XLMBL3CAzIdBklqINSz2/klFmYrFZArA
1JJe1GIIq+zrE1AUBEeQLKWwzA41MtXRnZ0B+IjEH7R7sEx6TNQUH5XaHCMKwmcGzIcfPzu1G2CW
4r7XPFBoonC0iUnBJ4syPxAb1caXw2UidDw9/jDs8dyOtv/+jEqz6Mwhtde5dkd4hDfwdRymNlCb
XJmztyflVX43H0LGMIjCbBE9NMmz4ZLyvFhmtKNr5E8Q14CS5p/kbFnZJrwWhprNduN+i29k+yVt
ZbwpMR/zpSOGqm9YSLGd+bHKjj89GElpkYsZipqY//wMiQ+8QpqghHIkzRap6J5s2SJ9Bb/cew1S
tFsRlJyt8nDXy12bvkxWfUFxgsnEYkjvTI9CZIuK70WGP2gFjL32CTcPmhs/5hvRuW5PyrlhtCg5
twaIikrWYHVpQ0D5cGPmVzdvUGKNTITnl7O4M1Z0NbMfd31tNHfSm5ONbjBZiGsAWtnCxqRmOGDp
90EYdeRe0KbjYMHk2YphwgjX4YSy7dkyQ8BOmX9AYP8E2t7pJVMtXAC/raI+aH6CPsupg9uaDJYY
ni5q/eTj2lCvIDChXDotPa8S1uySMlLkGyojVRHM6A6RT6XB0UjsmCawAEUDomsaleeuNXP0u+3l
i+HHXSTmIyny+b/ylfBg10kVVkXYDpAGlgx8PhG6QHz7SmBPSvZoJIXwDUc2II5Sw4WGJSA0mgCm
Hr1FBDTV2wgmdZ48695Nm1gbk+bFVxkelS40P8vTetWD+YODalJbx3lmMslfWCRPYqr7RRRdU0j+
Zs7fIRc0WMIcCaKEvJjDgYt8ajfFPtKqZjX1eHQvOJrlfPX4NzJLZNgW9S56WtuojUB01Omif4xY
Jkgq0VX1bnatAIFGuVlr4AL4v3tMAIIuUK/ynM8uUFJ+4wVjv2UfCemYL/i/DmdFAr8nJUuJCL/M
HsNplpGzpJl/e9Bf4t8zSPnGpUagqqLFKlFOAZ7MsakhSJRu5hc9rTAkuFDJGCqFnJC6zQt3Xo6c
9Jr5CJ8cdxp0GtIGxrm3STNCo58XlOavLssYdiCRGBkWEb5sukNoEWlmU/9WjvadRdA1gv7j7Kh7
mnHIGOJx7RMZVnRHUvYbUG9jlu/LTMKMhaWK3bjfji6TvC9xUCdZcvdDCY67IchBL73Vzn/gc1au
nWll7cP0IGeKLFBkbazssj4Mgh6XZ3z2CPIGg8Rj4p+/R7VuV2eHWxGKWoPYYzK6VXBSDdFSJYPF
+gjc6xdMf03tw7Ztecd5XUHdUy3l8ZG899U/g52dMzbuUdY2qcCDA8YzXDB7AdY3iwsqC6rr4ae8
PpRZaDCGkGPkhIZ9J8GLfAWsJXwBsvzjH4oG3kskMAKHH4C2kV5NAjHvy52aap+t7Bts2MDdIXqb
n2d8CwtLJ2pWh5bkAcusnNgyv85DUtlcg+VW24kYnCToSJ1qe+5vJqLYBYa2BIZnhCGwJ7eqZPJH
M+o+Fd5MVhvrUDO9c8DhxlxbQA/EDpL73kejhrN7aW4ItF2SxqKaVGq1EBoLocNKpW2c/yNy+TTJ
gH096i3/PjGit4KjiraU5e0XEFEwI/cGjIiAvT4ymrzpTyQK0/rry+YT54beWSgqymuojOKTD2jx
QeZjone4Sp2PgKqH3kd7s50xH6B8tYsSz0jrAHiLlWAypY4PLLskAGVyb09i5OErULTbNd+wmSvP
OGkG6qeDBdmIGoQzbdFLqRy9xB/NMmoDyttBzVr645c+0XBxFS5lZCbejQPXiJ2P9OpWGtZtzWcH
wuhYQcXNe0Ku0lHCnlzER8OuS/7G8+Ld5xrvybuAPxMggbi+Kos8+VVHwRCk0O3wKsZ1afOpEYw4
SjQQNLFjtmmIdL+GuiLKWDjYoeWdcQPnTKQ+r/Ry/h5Z02k8CEr3lmR8cAiT6xWDQDZ289HLB18D
v1LgogKQFxn8jlPTlXkMxrgg7+8y13OHOfE5arPpIsVwCJunyZiuqZMeDLvF17nDEy9tg48w7y3f
f4y281/Hn/QzLct/FHZgR5snIEc5jpSPSTAoQ1SsyW/8FTHj0P66Tr3N35gyIbijjgCkZsi03cKb
9WOJlHgGH+K5DMFSJpqJxMsGwXcW3TKah9yJOdvhqL9F6RibldBkM1V9d/UmGXPDzxqBvZz7iPEi
VvqCpkyU+joSzKzaodiNtgkgk2youONunJOR/cky0hIXo3gMHhFIRb4ujq9BBjoPN1Lht59ene1r
g/26n1u2FeBbjL8HiuJVIfRgfE47Fuc0xvM50nw4v8Fl7XgNJYW/a5Vb6HDATnL6ykYgtZcOPyo3
JPiBa0aOcBiusuvL8rIIYXrUReylviDQTcU87vJ3E4yFNBn3EJldEMPaMNnRjJ1WNGjq0Xd6uo7h
YgEBbnyVlwP8TbY74GsB9uD7G4HCydcKQresJZnqMv4jnDnD66+APPnYaQmQN7L5cxM1V/pARe5y
Dc6C7S36+OyPyhKlkhDixY8GEywq4Mp2cEE2gKWa0O38eCZ0tb36/Kw9nw0QPO0tc9xVM4K5aKBk
exI/xnYFpy0Y29zESYM+JLC1mFdx+SdSy4wLaiP3Z+3sBhDTfTn6MDEgJ1N5uWNaYnwvg5ytu0A8
mGuMfex0/zfVDGrANkFbhKFjsLNKtURE8y7aC7kJc8k9ajTeIXWYL6x9QpoJmriHsAWb6a09n1yv
RsDtrWXnsdjgYwwcrDTu3b7wtTaSD+NKQm3HfW+JUjsCC+1ODO9EAPin/pIJoQy5lMLN1E7950o0
HKvdYeNtnJUIEVLB+STGdrFBV+dRpvaKYY6QmtAyvosnym1Az8HRFrZ7y/4hQX2wLxiyG9SlWCfJ
UnOUsQyTuGsR6O5fVMap+ekXEwO/98gn74iAzxpm/cRtdCL80q/FEG3pz+nylEeOa9kuR0a/l0B+
6X2AzU/zygIvm8H+klRLbi5aUExAVjVBPFSUoP01cYj5aZeSIRZR0ohw2hMATd2aJU+2UvHks9wq
hMrR+XjdAOWNU3BZQdUYVBtG2V4IC4wLlSqaFucdkNAHs2XJWaOiqbDizHv8umcVkVLG9zr3QAxY
ntoEDw3Bjblc2VUtld2NzJ2+fw5EsxmnrqRL40lsFHWbjvYbqqzwJZPLaNikL6HV/QOvHc37Ezu7
Ja2VOLFc35IaWIr6YB2k6K/Xo4Bs4Nbztd8lQldm8ey4FWtkRur1b6H7ED3A3qTWmHjXgHFNPQTY
Rz/4EVCZSMV+hscRGspCAN/TIlWeSsOBM9UzE6sANOjR+f6Rl/ngJLCCdglbSHWNRKhInxo2fgPQ
aSpzt3qcUBnfVGN37tS/Wzr7qwDlos98Q1y47aRtSb17I7RNBTKHvXEcfsBO5Yex9fMuF/PUXics
DHnP9k0CQb+ECbt5+7woXN6d76Z49aGvZZLONwJnE3GL6H7uAmLXp6enRrOuIFtxg4uBYBd31cVC
sLZvbaYTZKsZSmlKSiqjH+5PNh6WFixlveEI5agTPZPV8ySFjpuMdBLIyuZJ20yXccWggktzozkF
17BzBNSwgpOGvFTMNvYNQKS6oaCOUsDGGV0pcNZfTWXvFoAtVciLFy/IMlSb65x2K9Co1x6HxkAV
IvpKQOOBPQWAhMB0FPsd6wSYItbjOrufJZU/deGWHASpy0L8WxURa4bvIHG0bkYcybNdcqywAMxZ
uX7NFirt3WLnXQWseU84nAz7uGfCpBWe6ztwNLXt47Y4XbcHvqYZRlqNB8FDluhvmO7Hj07O+gqF
i5XuRpvEgK32fwgrUFIFf24gCQbhxz1VxjFqI+VjEmyGV2RXbEMP0CFTKphKEK96Kle2S4AduVnU
8XW8tZtmsvOGrEFfQ/aPlp9iRX+V8++WGcPMFSpPQUxgHfxm5NrtO5taO7JyWdzq2Vp6QrvpxgLF
IZe8M/7RIbltl+vDapNs+oBpBYVysyB1CuEm2CI0ApZp3k9uCRwdfgmfJTC/0L5vmmUEiI8pA84i
K/nUCiyy1pJGKlK6DCMd+3FsR5BwUkbk6TTp5KK3nQ14Cqn6lsaCpY1D9KjxOu69TMIhPm9qzKLY
k1mwNUG4kgJyIrOZw7t1Ngma4/n2MmW6yDsQCpBM4fUo8LRtFJ9d7fvvlWNdGEnIw5g+A64hZS+p
ib7lHHMD2vQwZlw9dWsSZXKQb1g66gWeBOni+P/jVnYcYM4MFZ2DivJOTTqAnRjyIAGOH/D792tR
4A/8fgbtmxZfNbw/Z37w+9Gr7ewFT1U7dvORLKq+MtLELN/sF/ZszwxKCpcYfGObWEJUIyxHQC2R
lgctrZ01CY4WwaDzCyIZ7Y2GuJJ0I2lPVvLZYTs2MnrMt5hQbTd9pvehYOeYI9gQIB4s3pwJ8wZ6
6tQ3YsqPhwzBHb817LAqHXuNgb7+rUmVV2KPzqBXw6hXwpj1Tw7RUOfLUIBaO2yB6v6DEkehiAiv
KTSqChOTfV4bRziYwQsyieiUdQiT2faZI4n9t9iFmsMa5MKzABaIUc9Yn169pFb3Cb2j5WLqa3Sa
r7shIR3+4okousBRF93x/GEXy2Urpx5bwNOlluAdNQXnCQuF4lEHrz6rJvem5oA/LRwDhfrYQjO+
Bhu+4aU9tLBLTL6OuJlgYALtBYm5VR+SUtpyfUcP2alduJV4GYRt8ahNKGjskbqs7jliczACtaX1
KC8CtKHC+qbJ7F8/Z8UII+YUsbDJTCV4SC2b1s6CtTa3KE63J3vCDTI1AwPmqIeWPU7QoQ1lWG5V
2NTEOJG60HixCksyVZYY9q0BTKJg9sqmjylGKnRG5SbrBlM7XI9UY025W6EJh6p6eIpLqgblCKwB
SFa1jCQbFt4eYCq4V+vJf3zF+W5NlCoGlTO7g+hcQsnZp0E9lwwhgi6NeLPaR+ZpaCrVZHLddDYm
5RZ3y/QavW3Lh2A3sJ4MiEdaI3Nic3IzMnlfw7tqocJbg1NtjxC6cPn1tBieNM4i5ERZZQ3OpljH
c20YPuQ3/ZsMD9G2jYwuT+ltiWt12/uV8sTajuzivF466SGaMX40AUhhV99iX/KzpN7Cj25sgPXQ
1fKyh/OXKblmXJxqYP9y41tZwdDs5pTezmbbvLJozHlt+e+Hs9ZkbyLBE+99nc/4arXrPmiCTyA8
BBBBrCnl+0t+iluIKFNrG8nwi6b1hsqRdwMblOH0RzVT1h4+Nl3e/15iEkBjxo8pDlakw+rQmADU
2b9RyAjRM/EnMXCQAGhW5M9sxAv+3N122V4zihiPJfh6HQE2vORkO47KfbwlMTvrZmpGSo4nCTVX
I89pl3ubj2wN5eDBXoulsv9rIOZCWimMHUlD432ZvhZvbTaVR+cWS8r8Do/xpSV4YqMp1zkL5QdJ
7cnpAjbIv85e1cxqnBmnUaWvqACQTqcrhOgdabccHzDBsHlmV/WU6KC9VzKBGttny6UoPz2bDUxa
lXLqkscG66hfmsJ+FmClzuSDQSwYxsDs8MGgu/l3HDG+btQN6MD0YDtKwn0+mGwoOCh4iyA+boR4
ffxf9WKmMtrnNVQtLdjYfl1ovu0ukYDlunnu7JmAAyeDlBEx7fyuxoLVEtRW8hsV7KLRcmdDYn65
MUtyi/h/LcofezlCpX7YcimAcR8+heQnJgs5t/x6btkOGqnCQ4gA9MKlLamlglLL4Fviw1t7jcw7
QZrMtZxpbnq8CjRuotKHh7piYedN/wT8s2dkD5kjqlptaJpVpvcxTxC2KCqEWoI1HM7P20Nj1Xrb
3fKf99yO6vM1NoyEM4i4QOvWz6ZXaJi70ZB/jqWHd0JFA9Sr9N9vzjhChj3gAfRiPy38p5oXKs1l
wHU4CzddsP/DXghIk1F4Gd11kVyz4EzLJlhOzakze/GxCUuezV9YHgSU8qObBAaW+P3JCAwKP6Zj
hBDvFhgKeZ1PWtXFrz+TP8IbhTEVY8tmbT9ZYBl46OhkiXea7zJzQ3UrKsMWXz5DyUrVqRy/5O7H
BaC86prsCZrzFEdo+OGXlFTbmrsiyti6Cdy3hx7QMvqX3Dc1+WK9mweSLNwOhArpegYFpnJO7bCx
zLkIpp2HaItgH52LKehBUScfo5Ld+h/sur8rlkASfOjlyWcpnTXuvUq0vqC6ogwk3nKs7V4lkene
ECAAl7N5gNIWbpVkyNfHX+z0j8XCKiimRM7zPSLl8M97sXr6YTRda5FL/5UUlcXvWYbcCBcVldki
2wzVtOmtBy3ETBeM59Q4auRDbQlc4V6+nuWSSHV9YvwAErXfMVo4UXKZ8cs3UeD2AJBoAjw2msbO
/Yscn42NZPzOphiJf5ZDNq4WCG6cKqt2228Dt9e9uk0V3xgz2PzSA4mVjybEZYrx688aJeeT0n8Q
URmYrmphMc5zZ5hHqvWHD5NsKbOpd0ayXExrU339C2xjeIPgisXqzcEYERtFH4vk3xynOKJcLi06
fe3OPFhIcvmFo26PaonWOpEv6uPulFxRI7vTeUDzN3cwtYHn7/R/weM+MBlw938YTeQZRxq9zMD2
HStKNG5da4E6RnmBcWPwrNGltukAKCyGRXQp8DwAw2nAUwVPvs4zLqSjFHR5hdkq0+VbJsCY79jd
Ps1BNwNqc4Qdr/wowXqXCpTSpcSdgKiQ427YTTTkYAoL33FyoWvofMTkT4j2bQVkL7Agyh2yPKWs
6WOx9pfiVPFcmiK9tOtdYT5IG0JYkZhFPs7zDqIdecwjUZHLsVGc3xFUv9KKMpASF7QjecN0WchB
guuIghAXE1TX4oQCvDLQJeCyx8tvBiYUzsMe7FoXPrsUlzn//n1gUBjtrTGCz53z5/aAVNZoI5WG
jskZKi2ccEPqwprbPuXuUS1MkNexNLTIOE4qMOxCusmccSA8zK0GA/76lYNTXWSZEPQnoWFLOUyG
sKgjqP2nS3yRWV0uGrA6SjQQ7tf4QtEDTwu/5tfrmuGPnH1kJvclJIu0zx2HHdYO4Lza1gqkw/Dn
ARzxGqmAlyK+GLRptHwU5L7+5UvqDUs6sIrFl3RrRY2Yc+2hcslt4c+bdN5Sy69RBWF3X2LctgpZ
vPWSt5ioB4qESofg5RCRWvOqM6Uod6Ik1f+B+5nYKtUHySoqOe/qXI3cZBVp2TiG7pFSzTdZ3IlJ
pji9Ucmh7uIedsMQUwbQnsbD+ILWqntfH0HlHzdk3Z+su6rhx9rDYZYRYGqnb3+K+qfaZNX8YwGL
bTxWfUkqS2V65cRN2PV1b+EjADGy7XYF/m6bmC2pK+mpZzqJ++Q8D+VT8FkCb2KsvvbOIxzATvtE
YD0iKdJ2xwizFxP2+srtUxrQN2kuCu515tccQLvjsPAAqaPW7AfKEN3Eri5vQNiHbL0iQ+PR3bh9
uRo0KTXBzB80Yru/QmUwpLb3RouapIcFBA+n0F2kBIQVqmcnK123Ckw4lAAjr029SRePa+zUaGV2
y0868kfNsOwmtVYyXReVrFJ3xpLZwa6OXCDfo/H/P0dDB6zgfPDA2TEzyGKb+hNlf+9ElGwowQyW
yfwiVMW2b0N4wQm+S1MChUlYV2uAEzi/oc8kCS1BH2MlnJrX/jMK5aH08FfbbGtlkabUkxyp9n9B
REYmqMRHxDzoqoQbYxvfchYYaoGTI7kALitslv4bWFxVCKwVDbbOYfs09z1GxVGsPJgeJWsKxoRT
DTtk2i7qAH/1uADYQ3ilUvWshoj9ECpCE0nIkFn3NQ6K/8PM68qxQGXwqBEPvH2e6qA6l9Cohvkv
Evub9z5kKD2lLeR5Xyg4nervvtzrdoNyXFIf/ZuUF3UuamdPVcz1qE7Kfwgdurrejh6qX9cKYoPA
WHKNpv1T5FDIfXxPk0Q1tocCLhtrkjV1VuzZHP3Pf8NQowl0sUw0tXZ1h2ZQ/S1HJiGwvg3FOevP
+Xt+8hnH3g+SYmmiAz+psGZScIKWC8eek6hHONipd63ds7chxpXAAzt5ONDEGTmG+USWzQCXuq2v
gDkw0avIx1l0CdIHgu5Q72vpOOXBj0JBWKwp5f74ULxMS0IA6SfIGfhwoqN+Z94A6P/FSkIG87zf
2DskqttbXvFeOrdlP+nVZByESPq2eo2WoqqWonh9QAIh542z3WW6ITggBRxoftORSw5Qw+SWISy3
AdE8VH3E381M1BxjGGEV85reLeBIHOz/4VftaZGAUv0xmIsp7vtmsgy94LzDERAyCba0EbSXY/xn
tQ5h3OZaLu90n4mmDzWHCGXo/JSQjJPrfl2lU+FFGuDN2Y5XJCI289ZyJj1zlWhHPCla0AvYDBIp
mGP4Xm70+/H6XpD79oOJejKXxnqeTrGTkl+pPKutciy8ShDVzyQ9XgwdxVYSXtXxRH3vkBt0ztKK
kKF6tQz8bVwjt6FQRsyFuEHaRt2LbzKtRKrbg312fuF8qFGh4vo39cDdOt26hA1ifv3HOEXFOYSM
8Ua/CBiLPqgIqf4M/sq4JV5L/VMdTbl1qm7rmm+lInoolAiaYKBplhafV86HVn2rmQVB4B2ABhn9
6hhP0qxwH5T0bwvMhkQpZvA6IrYQH8qKEMZt3HfCb88NudE/fQ58O0ai9oOZPRbZmjSrxMSMKvi0
yKPy9jaEfqKtvzOn6sO38EOzwV1RiuJ3UvxgaQphps7/i+w+9ZwWSeU8h+Yi0yehq+FmP/iADDYL
zkL1ZOFrUB3FuFtAN2NiUPNkqMhtYZEdUGzA76h2EA3BC1RxFEaQUlEYZfD0Nkh23F58eMLpTsLX
Ea9Lwl0m0FLoV6fB7f2gCzaKEABaaSDI67QCyID9/hocaTKsWIsHDIWdQEUMKKvCr41OtH0cphxo
sEfgfzf4quS5pMFy7/iqWyCDEY+Pg9mjo/Dta8aBHdG48hK0IUC6RhyJlBQT8DdvsBBwwosp+it0
4lil1VE4Bw5puWqdpg7ri6fhBEZx4FzxCbkohE4L2PyDyzCWTPsJJeXZ/AlFX+1NVF9Fv2+t1vzR
S/Kqw51m8Yt3D5n/qblqf7E/431lFeUzrcIb7t3f0xB74AdZ7xFjEmHLSwp/+p94VdvL9rQQW0Gf
+4llryXSBw7kjwYadPYcFATBA0B4bE1F3MSIzt/Pcsz6MGc8Vgan2nfnkYsWXQxnWMfHRdn8YzJ5
WIawv6c5E+BWpDnRu4BY9xioFtFp9e/4tCX8YBCT6ih+SNiUwPOsGEE32vYVqW6CdNNnt4hbuyYf
5Z+HQCvRXFRv3mM9qTZ/sfRXFV1jehTBYbd8NbD4mLVHx9otpopsPQmrSXDaQWNA0gNgqFSp7Ck7
gyQHV2e19K+VHZhd/1Va4D+eTwOu5NIo2gH+qKdlDPAO0N7M59QbUxsAtLPnDMR9ymv2KNS83Dex
oR9m8l3tFqDz1o7iONYkl4tRKDubWJQj5m+47gwgmFjUwD7dJSJEJ8aVR0dTThkiGnrjqQ0cjVPI
LF1FWwWwFuK75r2NXkaU662ZWsa/ZlhY5lbrvwL7P8mPlNNsN7EaX+uJ0ScMYcPFlVElnk/lgVYw
0HSvNe45h3aKLrllpjeOa/X8mnx8C7uXVmLV8BII36IbbodjCpvWA7BJcaJmJvVKF9Up6OISqyPd
TDKrkxACWaxxMFjsUz6gx9DSUvqzFfY+zYLavSjbk/sIN4sQJ55F77DzNJpL0+xxCvYvhsoQzoj7
a7iE/1KhAwHCbbm8hoP3mDzNpp3ANhPpbCeGP5dzcU/pzvAMgpRUBnc7ncMZ7ySTIhzEQXAeKaFk
Dfqs3pHeyvNKn2r8v0d6vCk+GDDUoI/d6qXh9tKqiy+TALMXNu6H0IT9wl2hsikpyALMOQ4r4v1E
fjhCcsT1HSdxgDJVvpxOcXZcplH2EnfMbRcmfgeTDkh+TOiTBj7wIkCWJhI2WLT0Ek81CX3vVNF7
9HTJUNce2PKOUomDVUp/F09+yPQgfqv1zHcYd6MeTgyxRM2qyl3iNwC7STxqQwZp+DHLpGmnEhGr
valLrTZ/4FIkOy9e4ckxPd78Anntpf0rvl3SgwnWoK1uJtkVpEYgiEpGrvXX6YeOnQHTMDe7C2gH
HmnsqmHumcXUAjsajrJ2kg7LwKQgmwKItjiF/P9q/XiMYDmx+7pudXnIx2pB01UrKtiZxZNRlICv
rIcj2K+6yqNLTaK0TSl8PvHbqQK8caSb8HHdBSG5a9wR+05WhI4bzcSMiU99yMae5igd5Bpo1+N4
9h2nI87nbnvStE7qrfqsyjLSA6VrPZYZDxxfdM1rTD/ly43ZCeB9K4VgXj0NuwaZA1b9lu47kzgc
UULBJey2/oCM52ax18kSYQpm7gOV/iHSwSZuiEok5FWfarLcO+aow1zwCsMp9247enV5wAD045sv
WJ/6qIr5qBsXvOQw9LqctPjKXSTJQI0ooGqk7qBxvvF7kvyVUyvK5yWsJqpKYPZ7u5jx8hRgxeiJ
9o1TTCQd8ZcWubIzt47UkbruHjeECJv2JHbgtB9WC79aMmub4Ol/PGxYVQXxu17KZLrM1jzhSUL+
AXre7V5z2BIDE1n+hapqykftNf6PYpsS04BoP5nHCJBGuONWX8eY5d61lyjsxEYo8mgZNSUP/asZ
KvAgDLj45yJbNSK9HMr00arW5UHN1EX8VxJDqV89bJAxvt1e/XdYQL7dwG8hRL42Bs9mQrGD7QD6
DzK61XqquCZ+/RZGqob9YHWOnCem511kkdWUrQzgcLMO28fKbSNeQmWEjjCy/hpID/wOjDHaBq78
4wbY8ZhG6qmvSA+uUfyxe8s1cr9UkRCHpSj96ledt78WTAGiIsM8CvH2WLDnDXMFlzmCI3T25qD+
j15KMj1g3/WP24Yv8FL6TgMCeiXvnTeCQuxbYeZsPYi4ITsQi8S8uuPr7LwY0qG/s5jU9B0E9Miq
uWmlARvBWKD1uJqXhtMdjFxtaodqp/vJxXfAmIMw7Ykmx2JYe8BJNRfSGUyuu7CKNjf2hy8OTlKS
S6JbupIomXC7H+w8DDP1CkVXvcaKg/Y1RMgeOU1MtPYxaHEqouQgXBhMu32phB3oSBYkIpA+9lGo
SpuS9g+Rch316UnkGK1qRzjWKLWGsW+YQjTg+zkFQYlxTGx4F6KeGMUGM/I9tKaAygXO4jpTpyjM
7KefZL6hJAi5/DxsDM0oWTvH6LVa+w3V2lkqI3s6gHDC9sq49ERRG6TmIssGzPWCAqFER5E1SFox
7YfyKwc26rkvfZXPkLPdQbO8Nv8SRjJjBSCT+5UiLdCi8nHSSB8EcUx85iPbb3eRqG4JCr/Wpaak
9A8DDt++X7t3hVjQLsrYOJmhSWR106iYYJmFZ59jcUR0N7YwzvdS+EwNtcYngE1e1wWKCjuH02bK
KH9nJLlfZ/xjiVILuMEC0MFPkpnMwPVwhXwylo07LrmjwTbMiXtXAh81FsHj25PdTyQPc1x8Ge1e
mzypZmuEccZEJK/Ti49mOSboEy5Iar0fTg8lzQLxWPMeohsD1WH2qvsdfErqnpxwsgIVdhTKx+PU
kxpA0A6y0Sd/PwBmJ7kioVusYgDhl9aCHeD1BmvfhB3m3qnSkBe2JWz2lEqVd12FAljUbeaH0lb+
LnTi/19zGOvoNdoopLHhl+0wixJSa4Pni+lQsJdf07fHchHPHsCOkRTpwWctNz94gxfNfcJ2RCuP
oB7LjL770H3OA+vUu7yEi/hzAzOizd7+YNwPHPIJGNYhWZAv5oJsI61/kqIcMW+ytksX/+dJz001
iXnW1zlnSbgFdXsI+nZ2NXKP34NLcj5Az/PN31v5y3HqkmiWOxij+yuH82C9cJR/d/8z/pG7Vk98
7aXfvyOcxE8aOJturJIau6fJDW3sKOwrgfdEm051wsQdMzozZlIQx4FkxK+43RG51L8UI0rrHe9P
iAZ/rcM2F+9uB+nrbyBhLwf2O299ZlD3CiO97bivVuvO0dZPUhL0INVEy7aNuodpYuHF8LV9zKMl
ndK19bwwONNdEJB9D9JcQv9aIzUIiHthRC9rdFOwz6d2GntBByTM3IIrMcyNtGhl9tTkcpj9Cpki
9dKfQ8XbQRCG2B2caejmL7Fj22RBj7EGg2Lg7kMQiqNaznQviC24tKQsTWNWsaFBViAquVsVuAL2
Jb72OFsaaUGFMb3h19zcxdKmOwypQleO/vLZ/448by9135G/h0fUzdIc01ZPMZ7+b9EDQgoC33Fm
K8kgKCXADN5lLzrKr1h9IxhcqwvsXIJGRs2xGcq/TvAgo7Pvk70ORaWSf/b6aUCntXZmNwB7yhaM
1woBzMPhF4AJDCvlpl+nALQwLt5oHMC20bl9GdmpBByhkyd2SwGLXJxQj1BIsH75QEnD3JpezcPi
1XW3uLT/OLOhVQFMY5upTEylRJx0e2aQb6w1EERjhdNOtYqYSQLOUszbyIYYAeDmMPcKx/dpT+3X
56rK0qb/s+WjLlxHPyoYTK/nUX8sP1mAyyX2f/Xm249RHKubb0L8mMakKXQ59JMQ68Z649dpdDQz
m3R36YYOXYyNZQ+yUr9/y5T2YGhkks7HKHMr4KGKUoK+yjGoLucQan2kucn2Ajj+kAq5GMy9s2EW
D7tsZ84Hvh8CWh3oOz9EYpyjVjsm0MgK/MQd9E7Qo1LDw57XcFZcmO87iIY0Rey7UuV5vqpxwz3j
I08vByoQky1CE+mMiJki7G4hBcNdkBlJtzk3p24DhnvUlGun7HuI/ZyZPyxb0+/MOGXV+zlL8EDN
tk6sP4Q0zKs/zO6eSTPTmmfV/6UXr63gILSSpBKYG3NdGBAILICCVrvtMEYP7rkCVT86tpuiNYY9
x5dACOq8Cx7s63Zer/wxpE0DYxo/hzcFunEPx/HrG8Bj7RU6PfOo0W+tBElC9kgUhSldA15u2mX6
DVeHZeMg4O56L5uPQUFe2AREMWdJPUKmWPcg9S53vJFzjHTxyd8WZ+Cs4/dF3F3+LRwULURJ9oWT
5pVyrcEAgMwIWp2K7FlXOAz1A5FDYIL295nQHK2C52VDskWxFWYPw/N19s2pEeNjhJb3Kx6UeEUp
blNVCyMW6enP0XWG5ZN8e05XKDF/DlCyfVZCLp6C3elx10G6othNs7FDUfqe61/QhUpZN/44mLST
kvz0xaAy3VzAZ5mHX92J+s3kaf2AAkViesyZfZR9vY2SAykeertLPhBvbnjcapJwoUYsEsO4JPFW
TUjar85mMDLovCHl9e3GMES1RMRYRWqq7H/lFI1TGS7i2HrxjYBQ1/4Xiw938FUWkn8DXddyXqQe
ElT1YRfCxiyaDHxUhIIImB7APJOko5e438eQYWWhGnu9DUBOXQUOutWP4I2KHT+UHD1vy1KRrK6X
b2y3xOBSDimE6f4c5gfjS1GOqad2jFp0BCvxr8xDli6kwn20AmMMXMCKj9B84syDIzdcIbhuYUla
SHfOBQLyZQY17DWKhjXmtldcfw2rHCRFh+Cc5D2hA0QBaZtcoNneha3WaNi4CugeHSdMCzkeFI2X
Ke4E9guvLmjN6cCdDX6r3vACpolJUCJz8ZjshtLrvJ8AsO/6oaOA4PcDqozeBEVahz6h3BJbAKVF
cS/FOYUk+UrqvlRO6kG4YhH+a6BmCnqh7RLpoEzanReRiaAcqXJf2Ec+gWSBhOXVgTUxBok4hVDg
+2XfJfvqbnOQ8APTnzJAaenDWwU8VllkemleptiKMidN03XCvYjc0VijPqaiUaKleXV0qkSAAT9N
66GCx6qDde1uonXrJWlL/lK825mJYNVfKrpxIKpGSD0Tj326nWPnA118epGuUCS9dyY4L0uUtO0o
LqGQx7MJI6g978jBXIObjyCYE35jD6XZ6ce3gGurGchZNzLtCSRmJUwXorCrZBOTaqB8RJFFyDpJ
49l9KrGUhbqTQi2/GSeNSmnlx6EEB6uqMRu/pP3OH3fHmfREb2mo3ttI+DYA+wRq92EohKB2ePAO
7KE+pRlQfes5hkmpZGTYDNoNXNyV4IW68I1Jdr5pUlHWPscok9xTSPlHmAcxso4PQ6QBOW5B4l48
XaibBVscZR3WW3vY3aNxJQlrhsDz6KyOiwnmZXy9P3KIimkQoTryq090d420X5nm9PXYX7+7CD86
CJHTE2pR7puIhd7O3F9UrPiiuBLejwyfxCBdEifPKZ36P114DY7OjldUW/zrEUW41Z6mFfQw28im
AQR390OGphP8APUNJOk04EHMO+Z8bgxbV5QLlV+tEL5Mx7Eb18SHraYwoNMfq2MlnBK0h+YzRKK8
6EDccYAeYCYedyUPmTmkIXhyesA1//ydqHZCHbCe/B/m0r3rUYtvU23zLJd/RcQFKNPM/UFFLWCP
agsyNaGWWv4TNvT94p5pVe67bCn3d/0CvNULa8QoefhMf2ZqycQjnzspCwty9UO9FIee8qaiF61N
+EdDgYAefEPl2diOtWPeXeZkDK6nVl5qnfN3u8Nbox5NyL3gALO4Dxpqtft5sqPVtvulUuvKrABe
0Ok4ArcUL3Q/l9zB+y/WflIdjL3Q76TbkIhfo8oiefgX+66RH8bVHSPkwPpO3XlxVpmwmLu7JxTU
K3dIqnlWZ9Y6ukh/PKM3GusUfVCL7e+IYxE0DzwUJqoCSVO/bl+qcW13n9/YfbTz4ar6o+cdkU/Y
Kw8HdfeA8FDGpbYkZMk5W3BguLCNlpdjaB5WKPuD3p9iQoNwA0kZ8xDEhx+auFCGfB/JNfs+JNtd
H+h1Qv0hNow8V+8UlkZ6ki/bSGJLkyXIp/7HkppRbwSU41y8cqyA4TplRMMuRzJz6bo=
`protect end_protected
